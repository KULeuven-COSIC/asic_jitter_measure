* Top cell name: conf_128

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm5 net17 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm4 net18 in1 net17 vss n_mos l=60n w=360.0n m=1
    Mm3 out in0 net18 vss n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=60n w=360.0n m=1
    Mm2 net5 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm1 net16 in1 net5 vss n_mos l=60n w=360.0n m=1
    Mm0 out in0 net16 vss n_mos l=60n w=360.0n m=1
    Mm7 net32 rst vdd vdd p_mos l=60n w=480.0n m=1
    Mm6 out in2 net32 vdd p_mos l=60n w=480.0n m=1
    Mm5 out in1 net32 vdd p_mos l=60n w=480.0n m=1
    Mm4 out in0 net32 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=120.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT dff_st_ar_buf clk d q q' rst rst' vdd vss
    Xi0 clk d net17 net18 rst rst' vdd vss dff_st_ar
    Xi2 net17 q' vdd vss inv
    Xi1 net18 q vdd vss inv
.ENDS

.SUBCKT conf_2 clk in out<0> out<1> rst rst' vdd vss
    Xi1 clk out<0> out<1> net14 rst rst' vdd vss dff_st_ar_buf
    Xi0 clk in out<0> net13 rst rst' vdd vss dff_st_ar_buf
.ENDS

.SUBCKT conf_4 clk in out<0> out<1> out<2> out<3> rst rst' vdd vss
    Xi1 clk out<1> out<2> out<3> rst rst' vdd vss conf_2
    Xi0 clk in out<0> out<1> rst rst' vdd vss conf_2
.ENDS

.SUBCKT conf_8 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> rst rst' vdd vss
    Xi1 clk out<3> out<4> out<5> out<6> out<7> rst rst' vdd vss conf_4
    Xi0 clk in out<0> out<1> out<2> out<3> rst rst' vdd vss conf_4
.ENDS

.SUBCKT conf_16 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10>
                + out<11> out<12> out<13> out<14> out<15> rst rst' vdd vss
    Xi1 clk out<7> out<8> out<9> out<10> out<11> out<12> out<13> out<14> out<15> rst rst' vdd vss
        + conf_8
    Xi0 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> rst rst' vdd vss conf_8
.ENDS

.SUBCKT conf_32 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10>
                + out<11> out<12> out<13> out<14> out<15> out<16> out<17> out<18> out<19> out<20>
                + out<21> out<22> out<23> out<24> out<25> out<26> out<27> out<28> out<29> out<30>
                + out<31> rst rst' vdd vss
    Xi1 clk out<15> out<16> out<17> out<18> out<19> out<20> out<21> out<22> out<23> out<24> out<25>
        + out<26> out<27> out<28> out<29> out<30> out<31> rst rst' vdd vss conf_16
    Xi0 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11>
        + out<12> out<13> out<14> out<15> rst rst' vdd vss conf_16
.ENDS

.SUBCKT conf_64 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10>
                + out<11> out<12> out<13> out<14> out<15> out<16> out<17> out<18> out<19> out<20>
                + out<21> out<22> out<23> out<24> out<25> out<26> out<27> out<28> out<29> out<30>
                + out<31> out<32> out<33> out<34> out<35> out<36> out<37> out<38> out<39> out<40>
                + out<41> out<42> out<43> out<44> out<45> out<46> out<47> out<48> out<49> out<50>
                + out<51> out<52> out<53> out<54> out<55> out<56> out<57> out<58> out<59> out<60>
                + out<61> out<62> out<63> rst rst' vdd vss
    Xi1 clk out<31> out<32> out<33> out<34> out<35> out<36> out<37> out<38> out<39> out<40> out<41>
        + out<42> out<43> out<44> out<45> out<46> out<47> out<48> out<49> out<50> out<51> out<52>
        + out<53> out<54> out<55> out<56> out<57> out<58> out<59> out<60> out<61> out<62> out<63>
        + rst rst' vdd vss conf_32
    Xi0 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11>
        + out<12> out<13> out<14> out<15> out<16> out<17> out<18> out<19> out<20> out<21> out<22>
        + out<23> out<24> out<25> out<26> out<27> out<28> out<29> out<30> out<31> rst rst' vdd vss
        + conf_32
.ENDS

.SUBCKT conf_128 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9>
                 + out<10> out<11> out<12> out<13> out<14> out<15> out<16> out<17> out<18> out<19>
                 + out<20> out<21> out<22> out<23> out<24> out<25> out<26> out<27> out<28> out<29>
                 + out<30> out<31> out<32> out<33> out<34> out<35> out<36> out<37> out<38> out<39>
                 + out<40> out<41> out<42> out<43> out<44> out<45> out<46> out<47> out<48> out<49>
                 + out<50> out<51> out<52> out<53> out<54> out<55> out<56> out<57> out<58> out<59>
                 + out<60> out<61> out<62> out<63> out<64> out<65> out<66> out<67> out<68> out<69>
                 + out<70> out<71> out<72> out<73> out<74> out<75> out<76> out<77> out<78> out<79>
                 + out<80> out<81> out<82> out<83> out<84> out<85> out<86> out<87> out<88> out<89>
                 + out<90> out<91> out<92> out<93> out<94> out<95> out<96> out<97> out<98> out<99>
                 + out<100> out<101> out<102> out<103> out<104> out<105> out<106> out<107> out<108>
                 + out<109> out<110> out<111> out<112> out<113> out<114> out<115> out<116> out<117>
                 + out<118> out<119> out<120> out<121> out<122> out<123> out<124> out<125> out<126>
                 + out<127> rst rst' vdd vss
    Xi1 clk out<63> out<64> out<65> out<66> out<67> out<68> out<69> out<70> out<71> out<72> out<73>
        + out<74> out<75> out<76> out<77> out<78> out<79> out<80> out<81> out<82> out<83> out<84>
        + out<85> out<86> out<87> out<88> out<89> out<90> out<91> out<92> out<93> out<94> out<95>
        + out<96> out<97> out<98> out<99> out<100> out<101> out<102> out<103> out<104> out<105>
        + out<106> out<107> out<108> out<109> out<110> out<111> out<112> out<113> out<114> out<115>
        + out<116> out<117> out<118> out<119> out<120> out<121> out<122> out<123> out<124> out<125>
        + out<126> out<127> rst rst' vdd vss conf_64
    Xi0 clk in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11>
        + out<12> out<13> out<14> out<15> out<16> out<17> out<18> out<19> out<20> out<21> out<22>
        + out<23> out<24> out<25> out<26> out<27> out<28> out<29> out<30> out<31> out<32> out<33>
        + out<34> out<35> out<36> out<37> out<38> out<39> out<40> out<41> out<42> out<43> out<44>
        + out<45> out<46> out<47> out<48> out<49> out<50> out<51> out<52> out<53> out<54> out<55>
        + out<56> out<57> out<58> out<59> out<60> out<61> out<62> out<63> rst rst' vdd vss conf_64
.ENDS
