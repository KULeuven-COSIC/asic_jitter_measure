* Top cell name: mux4

.SUBCKT nand2 IN0 IN1 OUT VDD VSS
    Mm1 net13 IN1 VSS VSS n_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 net13 VSS n_mos l=60n w=240.0n m=1
    Mm3 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm2 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux2 IN0 IN1 OUT SEL VDD VSS
    Xi2 net16 net15 OUT VDD VSS nand2
    Xi1 SEL IN1 net15 VDD VSS nand2
    Xi0 IN0 net14 net16 VDD VSS nand2
    Mm0 net14 SEL VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 net14 SEL VSS VSS n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux4 IN<0> IN<1> IN<2> IN<3> OUT SEL<0> SEL<1> VDD VSS
    Xi2 net8 net7 OUT SEL<1> VDD VSS mux2
    Xi1 IN<2> IN<3> net7 SEL<0> VDD VSS mux2
    Xi0 IN<0> IN<1> net8 SEL<0> VDD VSS mux2
.ENDS
