* Top cell name: top_level

.SUBCKT esd_pdiode N P VSS
    Xd0 P N VSS VSS al=5u
.ENDS

.SUBCKT esd_ndiode N P
    Xd0 P N N N al=5u
.ENDS

.SUBCKT esd_signal_4x SIGNAL VDD_IO VSS_IO
    Xi4 VDD_IO SIGNAL VSS_IO esd_pdiode
    Xi3 VDD_IO SIGNAL VSS_IO esd_pdiode
    Xi2 VDD_IO SIGNAL VSS_IO esd_pdiode
    Xi0 VDD_IO SIGNAL VSS_IO esd_pdiode
    Xi7 SIGNAL VSS_IO esd_ndiode
    Xi6 SIGNAL VSS_IO esd_ndiode
    Xi5 SIGNAL VSS_IO esd_ndiode
    Xi1 SIGNAL VSS_IO esd_ndiode
.ENDS

.SUBCKT esd_pdiode_lt N P VSS
    Xd0 P N VSS VSS al=10u
.ENDS

.SUBCKT esd_ndiode_lt N P
    Xd0 P N N N al=10u
.ENDS

.SUBCKT esd_supply_3_1x_lt MID0 MID1 VDD VSS
    Xi3 MID1 VDD VSS esd_pdiode_lt
    Xi1 VSS MID0 VSS esd_pdiode_lt
    Xi0 MID0 MID1 VSS esd_pdiode_lt
    Xi2 VDD VSS esd_ndiode_lt
.ENDS

.SUBCKT esd_supply_3_4x_lt VDD VSS
    Xi3 MID0 MID1 VDD VSS esd_supply_3_1x_lt
    Xi2 MID0 MID1 VDD VSS esd_supply_3_1x_lt
    Xi1 MID0 MID1 VDD VSS esd_supply_3_1x_lt
    Xi0 MID0 MID1 VDD VSS esd_supply_3_1x_lt
.ENDS

.SUBCKT pad PAD VSS
    Xi0 PAD VSS lt=69.0u
.ENDS

.SUBCKT in_pad IN_PAD OUT VDD_CORE VDD_IO VSS
    Xi2 IN_PAD VDD_IO VSS esd_signal_4x
    Mm7 OUT OUT' VDD_CORE VDD_CORE p_mos l=60n w=400n m=8
    Mm1 OUT_B OUT' VDD_CORE VDD_CORE p_mos l=60n w=200n m=1
    Mm0 OUT' OUT_B VDD_CORE VDD_CORE p_mos l=60n w=200n m=1
    Mm4 IN_PAD' IN_PAD VSS VSS n_mos_io l=280.0n w=600n m=1
    Mm3 OUT_B IN_PAD' VSS VSS n_mos_io l=280.0n w=400n m=6
    Mm2 OUT' IN_PAD VSS VSS n_mos_io l=280.0n w=400n m=6
    Mm5 IN_PAD' IN_PAD VDD_IO VDD_IO p_mos_io l=280.0n w=600n m=1
    Mm6 OUT OUT' VSS VSS n_mos l=60n w=400n m=8
    Xi4 VDD_IO VSS esd_supply_3_4x_lt
    Xi5 IN_PAD VSS pad
.ENDS

.SUBCKT out_pad IN PAD_OUT VDD_CORE VDD_IO VSS
    Mm0 IN' IN VDD_CORE VDD_CORE p_mos l=60n w=120.0n m=1
    Mm1 IN' IN VSS VSS n_mos l=60n w=120.0n m=1
    Mm17 PAD_OUT net28 VSS VSS n_mos_io l=280.0n w=6.4u m=32
    Mm16 net28 net42 VSS VSS n_mos_io l=280.0n w=6.4u m=16
    Mm15 net42 net44 VSS VSS n_mos_io l=280.0n w=1.6u m=16
    Mm14 net44 net35 VSS VSS n_mos_io l=280.0n w=1.6u m=4
    Mm13 net35 net48 VSS VSS n_mos_io l=280.0n w=1.6u m=1
    Mm12 net48 DRIVER_IN VSS VSS n_mos_io l=280n w=400n m=1
    Mm3 DRIVER_IN IN' VSS VSS n_mos_io l=280.0n w=400n m=12
    Mm2 DRIVER_IN' IN VSS VSS n_mos_io l=280.0n w=400n m=12
    Mm11 PAD_OUT net28 VDD_IO VDD_IO p_mos_io l=280.0n w=6.4u m=32
    Mm10 net28 net42 VDD_IO VDD_IO p_mos_io l=280.0n w=6.4u m=16
    Mm9 net42 net44 VDD_IO VDD_IO p_mos_io l=280.0n w=1.6u m=16
    Mm8 net44 net35 VDD_IO VDD_IO p_mos_io l=280.0n w=1.6u m=4
    Mm7 net35 net48 VDD_IO VDD_IO p_mos_io l=280.0n w=1.6u m=1
    Mm6 net48 DRIVER_IN VDD_IO VDD_IO p_mos_io l=280n w=400n m=1
    Mm5 DRIVER_IN DRIVER_IN' VDD_IO VDD_IO p_mos_io l=280n w=400n m=1
    Mm4 DRIVER_IN' DRIVER_IN VDD_IO VDD_IO p_mos_io l=280n w=400n m=1
    Xi1 PAD_OUT VDD_IO VSS esd_signal_4x
    Xi3 VDD_IO VSS esd_supply_3_4x_lt
    Xi4 PAD_OUT VSS pad
.ENDS

.SUBCKT esd_supply_2_1x_lt MID VDD VSS
    Xi1 VSS MID VSS esd_pdiode_lt
    Xi0 MID VDD VSS esd_pdiode_lt
    Xi2 VDD VSS esd_ndiode_lt
.ENDS

.SUBCKT esd_supply_2_4x_lt VDD VSS
    Xi3 net5 VDD VSS esd_supply_2_1x_lt
    Xi2 net5 VDD VSS esd_supply_2_1x_lt
    Xi1 net5 VDD VSS esd_supply_2_1x_lt
    Xi0 net5 VDD VSS esd_supply_2_1x_lt
.ENDS

.SUBCKT vdd_pad VDD VDD_IO VSS
    Xi0 VDD VSS pad
    Xi1 VDD VSS esd_supply_2_4x_lt
    Xi2 VDD_IO VSS esd_supply_3_4x_lt
.ENDS

.SUBCKT vdd_core_pad VDD VDD_IO VSS
    Xi0 VDD VSS pad
    Xi1 VDD VSS esd_supply_2_4x_lt
    Xi2 VDD_IO VSS esd_supply_3_4x_lt
.ENDS

.SUBCKT vss_pad VDD_IO VSS
    Xi0 VSS VSS pad
    Xi1 VDD_IO VSS esd_supply_3_4x_lt
.ENDS

.SUBCKT vdd_io_pad VDD_IO VSS
    Xi0 VDD_IO VSS pad
    Xi1 VDD_IO VSS esd_supply_3_4x_lt
.ENDS

.SUBCKT padframe_v1 JIT_CONF_CLK JIT_CONF_CLK_PAD JIT_CONF_IN JIT_CONF_IN_PAD JIT_CONF_RST
                    + JIT_CONF_RST_PAD JIT_CORE_RST JIT_CORE_RST_PAD JIT_DC_CLK JIT_DC_CLK_PAD
                    + JIT_RO_ENABLE JIT_RO_ENABLE_PAD JIT_RO_OUT0 JIT_RO_OUT0_PAD JIT_RO_OUT1
                    + JIT_RO_OUT1_PAD JIT_SCAN_CLK JIT_SCAN_CLK_PAD JIT_SCAN_OUT JIT_SCAN_OUT_PAD
                    + JIT_SCAN_RST JIT_SCAN_RST_PAD JIT_SCAN_SER JIT_SCAN_SER_PAD JIT_VDD_CORE_PAD
                    + JIT_VDD_JIT0_PAD JIT_VDD_JIT1_PAD TRNG_CONF_CLK TRNG_CONF_CLK_PAD TRNG_CONF_IN
                    + TRNG_CONF_IN_PAD TRNG_CONF_RST TRNG_CONF_RST_PAD TRNG_CORE_RST
                    + TRNG_CORE_RST_PAD TRNG_DATA_OUT TRNG_DATA_OUT_PAD TRNG_DATA_READY
                    + TRNG_DATA_READY_PAD TRNG_EXT_CLK TRNG_EXT_CLK_PAD TRNG_RO_OUT TRNG_RO_OUT_PAD
                    + TRNG_SCAN_CLK TRNG_SCAN_CLK_PAD TRNG_SCAN_OUT TRNG_SCAN_OUT_PAD TRNG_SCAN_RST
                    + TRNG_SCAN_RST_PAD TRNG_SCAN_SER TRNG_SCAN_SER_PAD TRNG_SER_CLK
                    + TRNG_SER_CLK_PAD TRNG_VDD_CORE_PAD TRNG_VDD_DC_PAD TRNG_VDD_TDC_PAD VDD_IO_PAD
                    + VSS_PAD
    Xi19 JIT_SCAN_CLK_PAD JIT_SCAN_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi18 JIT_SCAN_SER_PAD JIT_SCAN_SER JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi17 JIT_CONF_RST_PAD JIT_CONF_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi16 JIT_CONF_CLK_PAD JIT_CONF_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi15 JIT_CONF_IN_PAD JIT_CONF_IN JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi14 JIT_SCAN_RST_PAD JIT_SCAN_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi13 TRNG_SCAN_SER_PAD TRNG_SCAN_SER JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi12 JIT_RO_ENABLE_PAD JIT_RO_ENABLE JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi11 JIT_DC_CLK_PAD JIT_DC_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi10 JIT_CORE_RST_PAD JIT_CORE_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi9 TRNG_SCAN_RST_PAD TRNG_SCAN_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi8 TRNG_SCAN_CLK_PAD TRNG_SCAN_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi7 TRNG_SER_CLK_PAD TRNG_SER_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi6 TRNG_EXT_CLK_PAD TRNG_EXT_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi5 TRNG_CORE_RST_PAD TRNG_CORE_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi4 TRNG_CONF_RST_PAD TRNG_CONF_RST JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi3 TRNG_CONF_CLK_PAD TRNG_CONF_CLK JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi0 TRNG_CONF_IN_PAD TRNG_CONF_IN JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD in_pad
    Xi26 JIT_SCAN_OUT JIT_SCAN_OUT_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi25 JIT_RO_OUT1 JIT_RO_OUT1_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi24 JIT_RO_OUT0 JIT_RO_OUT0_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi23 TRNG_DATA_READY TRNG_DATA_READY_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi22 TRNG_DATA_OUT TRNG_DATA_OUT_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi21 TRNG_RO_OUT TRNG_RO_OUT_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi20 TRNG_SCAN_OUT TRNG_SCAN_OUT_PAD JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD out_pad
    Xi31 JIT_VDD_JIT1_PAD VDD_IO_PAD VSS_PAD vdd_pad
    Xi30 JIT_VDD_JIT0_PAD VDD_IO_PAD VSS_PAD vdd_pad
    Xi29 TRNG_VDD_TDC_PAD VDD_IO_PAD VSS_PAD vdd_pad
    Xi28 TRNG_VDD_DC_PAD VDD_IO_PAD VSS_PAD vdd_pad
    Xi27 TRNG_VDD_CORE_PAD VDD_IO_PAD VSS_PAD vdd_pad
    Xi32 JIT_VDD_CORE_PAD VDD_IO_PAD VSS_PAD vdd_core_pad
    Xi37 VDD_IO_PAD VSS_PAD vss_pad
    Xi36 VDD_IO_PAD VSS_PAD vss_pad
    Xi35 VDD_IO_PAD VSS_PAD vss_pad
    Xi34 VDD_IO_PAD VSS_PAD vss_pad
    Xi33 VDD_IO_PAD VSS_PAD vss_pad
    Xi39 VDD_IO_PAD VSS_PAD vdd_io_pad
    Xi38 VDD_IO_PAD VSS_PAD vdd_io_pad
.ENDS

.SUBCKT nand2 IN0 IN1 OUT VDD VSS
    Mm1 net13 IN1 VSS VSS n_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 net13 VSS n_mos l=60n w=240.0n m=1
    Mm3 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm2 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux2 IN0 IN1 OUT SEL VDD VSS
    Xi2 net16 net15 OUT VDD VSS nand2
    Xi1 SEL IN1 net15 VDD VSS nand2
    Xi0 IN0 net14 net16 VDD VSS nand2
    Mm0 net14 SEL VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 net14 SEL VSS VSS n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux2_10x IN0<0> IN0<1> IN0<2> IN0<3> IN0<4> IN0<5> IN0<6> IN0<7> IN0<8> IN0<9> IN1<0> IN1<1>
                 + IN1<2> IN1<3> IN1<4> IN1<5> IN1<6> IN1<7> IN1<8> IN1<9> OUT<0> OUT<1> OUT<2>
                 + OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> SEL VDD VSS
    Xi0 IN0<0> IN1<0> OUT<0> SEL VDD VSS mux2
    Xi9 IN0<9> IN1<9> OUT<9> SEL VDD VSS mux2
    Xi8 IN0<8> IN1<8> OUT<8> SEL VDD VSS mux2
    Xi7 IN0<7> IN1<7> OUT<7> SEL VDD VSS mux2
    Xi6 IN0<6> IN1<6> OUT<6> SEL VDD VSS mux2
    Xi5 IN0<5> IN1<5> OUT<5> SEL VDD VSS mux2
    Xi4 IN0<4> IN1<4> OUT<4> SEL VDD VSS mux2
    Xi3 IN0<3> IN1<3> OUT<3> SEL VDD VSS mux2
    Xi2 IN0<2> IN1<2> OUT<2> SEL VDD VSS mux2
    Xi1 IN0<1> IN1<1> OUT<1> SEL VDD VSS mux2
.ENDS

.SUBCKT inv IN OUT VDD VSS
    Mm0 OUT IN VSS VSS n_mos l=60n w=120.0n m=1
    Mm1 OUT IN VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nor2 IN0 IN1 OUT VDD VSS
    Mm1 OUT IN1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm0 OUT IN0 VSS VSS n_mos l=60n w=120.0n m=1
    Mm3 net7 IN1 VDD VDD p_mos l=60n w=480.0n m=1
    Mm2 OUT IN0 net7 VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dec_stage CONF_RAND FF_IN FF_PREV OUT VDD VSS
    Xi0 FF_IN net3 VDD VSS inv
    Xi1 FF_PREV net3 net4 VDD VSS nor2
    Xi2 net4 CONF_RAND OUT VDD VSS nand2
.ENDS

.SUBCKT nand3 IN0 IN1 IN2 OUT VDD VSS
    Mm2 OUT IN2 VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
    Mm5 net17 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm4 net18 IN1 net17 VSS n_mos l=60n w=360.0n m=1
    Mm3 OUT IN0 net18 VSS n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT dec_6_conf_0 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5>
                     + FF_IN<0> FF_IN<1> FF_IN<2> FF_IN<3> FF_IN<4> FF_IN<5> RAND_OUT VDD VSS
    Xi23 CONF_DEC<5> FF_IN<5> FF_IN<4> STAGE<5> VDD VSS dec_stage
    Xi22 CONF_DEC<4> FF_IN<4> FF_IN<3> STAGE<4> VDD VSS dec_stage
    Xi21 CONF_DEC<3> FF_IN<3> FF_IN<2> STAGE<3> VDD VSS dec_stage
    Xi20 CONF_DEC<2> FF_IN<2> FF_IN<1> STAGE<2> VDD VSS dec_stage
    Xi19 CONF_DEC<1> FF_IN<1> FF_IN<0> STAGE<1> VDD VSS dec_stage
    Xi18 CONF_DEC<0> FF_IN<0> FF_IN<5> STAGE<0> VDD VSS dec_stage
    Xi25 STAGE<3> STAGE<4> STAGE<5> net023 VDD VSS nand3
    Xi24 STAGE<0> STAGE<1> STAGE<2> net026 VDD VSS nand3
    Xi26 net026 net023 RAND_OUT VDD VSS nor2
.ENDS

.SUBCKT nor3 IN0 IN1 IN2 OUT VDD VSS
    Mm2 OUT IN0 net6 VDD p_mos l=60n w=480.0n m=1
    Mm1 net6 IN1 net7 VDD p_mos l=60n w=480.0n m=1
    Mm0 net7 IN2 VDD VDD p_mos l=60n w=480.0n m=1
    Mm5 OUT IN2 VSS VSS n_mos l=60n w=120.0n m=1
    Mm4 OUT IN0 VSS VSS n_mos l=60n w=120.0n m=1
    Mm3 OUT IN1 VSS VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT nand3_r IN0 IN1 IN2 OUT RST VDD VSS
    Mm3 OUT RST VSS VSS n_mos l=60n w=360.0n m=1
    Mm2 net5 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm1 net16 IN1 net5 VSS n_mos l=60n w=360.0n m=1
    Mm0 OUT IN0 net16 VSS n_mos l=60n w=360.0n m=1
    Mm7 net32 RST VDD VDD p_mos l=60n w=480.0n m=1
    Mm6 OUT IN2 net32 VDD p_mos l=60n w=480.0n m=1
    Mm5 OUT IN1 net32 VDD p_mos l=60n w=480.0n m=1
    Mm4 OUT IN0 net32 VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT inv_wn IN OUT VDD VSS
    Mm0 OUT IN VSS VSS n_mos l=60n w=240.0n m=1
    Mm1 OUT IN VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT dff_st_ar_dh CLK Q Q' RST RST' VDD VSS
    Xi5 Q N1 Q' VDD VSS nand2
    Xi4 N0 Q' Q VDD VSS nand2
    Xi0 N3 N0 N2 VDD VSS nand2
    Xi1 CLK N2 RST' N0 VDD VSS nand3
    Xi2 CLK N0 N3 N1 RST VDD VSS nand3_r
    Xi6 N1 N3 VDD VSS inv_wn
.ENDS

.SUBCKT ff_ready FF0<0> FF0<1> FF0<2> FF1<0> FF1<1> FF1<2> FF_READY RST RST' VDD VSS
    Xi0 FF0<0> FF0<1> FF0<2> FF_NOR0 VDD VSS nor3
    Xi1 FF1<0> FF1<1> FF1<2> FF_NOR1 VDD VSS nor3
    Xi2 FF_NOR0 FF_NOR1 FF_NAND VDD VSS nand2
    Xi3 FF_NAND FF_READY net18 RST RST' VDD VSS dff_st_ar_dh
.ENDS

.SUBCKT dff_st_ar CLK D Q Q' RST RST' VDD VSS
    Xi5 Q N1 Q' VDD VSS nand2
    Xi4 N0 Q' Q VDD VSS nand2
    Xi3 N1 D N3 VDD VSS nand2
    Xi0 N3 N0 N2 VDD VSS nand2
    Xi1 CLK N2 RST' N0 VDD VSS nand3
    Xi2 CLK N0 N3 N1 RST VDD VSS nand3_r
.ENDS

.SUBCKT tff_st_ar CLK Q Q' RST RST' VDD VSS
    Xi0 CLK Q' Q Q' RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT asynccounter_8 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> Q' RST RST' VDD
                       + VSS
    Xi7 net4 OUT<4> net5 RST RST' VDD VSS tff_st_ar
    Xi6 net6 OUT<6> net7 RST RST' VDD VSS tff_st_ar
    Xi5 net7 OUT<7> Q' RST RST' VDD VSS tff_st_ar
    Xi4 net5 OUT<5> net6 RST RST' VDD VSS tff_st_ar
    Xi3 net2 OUT<2> net3 RST RST' VDD VSS tff_st_ar
    Xi2 net3 OUT<3> net4 RST RST' VDD VSS tff_st_ar
    Xi1 net1 OUT<1> net2 RST RST' VDD VSS tff_st_ar
    Xi0 CLK OUT<0> net1 RST RST' VDD VSS tff_st_ar
.ENDS

.SUBCKT nand4 IN0 IN1 IN2 IN3 OUT VDD VSS
    Mm3 OUT IN3 VDD VDD p_mos l=60n w=240.0n m=1
    Mm2 OUT IN2 VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
    Mm7 net21 IN3 VSS VSS n_mos l=60n w=480.0n m=1
    Mm6 net22 IN2 net21 VSS n_mos l=60n w=480.0n m=1
    Mm5 net23 IN1 net22 VSS n_mos l=60n w=480.0n m=1
    Mm4 OUT IN0 net23 VSS n_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT max_ready CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2> CONF_MAXCYCLES<3>
                  + CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> INT
                  + MAX_READY RST RST' VDD VSS
    Xi0 INT CNT<0> CNT<1> CNT<2> CNT<3> CNT<4> CNT<5> CNT<6> CNT<7> net020 RST RST' VDD VSS
        + asynccounter_8
    Xi8 CNT<7> CONF_MAXCYCLES<7> CNT_HIGH<7> VDD VSS nand2
    Xi7 CNT<6> CONF_MAXCYCLES<6> CNT_HIGH<6> VDD VSS nand2
    Xi6 CNT<5> CONF_MAXCYCLES<5> CNT_HIGH<5> VDD VSS nand2
    Xi5 CNT<4> CONF_MAXCYCLES<4> CNT_HIGH<4> VDD VSS nand2
    Xi4 CNT<3> CONF_MAXCYCLES<3> CNT_HIGH<3> VDD VSS nand2
    Xi3 CNT<2> CONF_MAXCYCLES<2> CNT_HIGH<2> VDD VSS nand2
    Xi2 CNT<1> CONF_MAXCYCLES<1> CNT_HIGH<1> VDD VSS nand2
    Xi1 CNT<0> CONF_MAXCYCLES<0> CNT_HIGH<0> VDD VSS nand2
    Xi10 CNT_HIGH<4> CNT_HIGH<5> CNT_HIGH<6> CNT_HIGH<7> net09 VDD VSS nand4
    Xi9 CNT_HIGH<0> CNT_HIGH<1> CNT_HIGH<2> CNT_HIGH<3> net010 VDD VSS nand4
    Xi11 net010 net09 net021 VDD VSS nor2
    Xi12 net021 READY VDD VSS inv
    Xi13 READY MAX_READY net018 RST RST' VDD VSS dff_st_ar_dh
.ENDS

.SUBCKT nor4 IN0 IN1 IN2 IN3 OUT VDD VSS
    Mm3 OUT IN0 net7 VDD p_mos l=60n w=480.0n m=1
    Mm2 net7 IN1 net6 VDD p_mos l=60n w=480.0n m=1
    Mm1 net6 IN2 net5 VDD p_mos l=60n w=480.0n m=1
    Mm0 net5 IN3 VDD VDD p_mos l=60n w=480.0n m=1
    Mm7 OUT IN3 VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 OUT IN2 VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 OUT IN0 VSS VSS n_mos l=60n w=120.0n m=1
    Mm4 OUT IN1 VSS VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT buffer IN OUT VDD VSS
    Mm1 OUT INT VSS VSS n_mos l=60n w=480.0n m=4
    Mm0 INT IN VSS VSS n_mos l=60n w=480.0n m=1
    Mm3 OUT INT VDD VDD p_mos l=60n w=480.0n m=4
    Mm2 INT IN VDD VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT wait_ready CLK CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
                   + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7>
                   + ENABLE_E2L INT RST RST' VDD VSS WAIT_READY
    Xi4 CLK_INT WAIT_CNT<0> WAIT_CNT<1> WAIT_CNT<2> WAIT_CNT<3> WAIT_CNT<4> WAIT_CNT<5> WAIT_CNT<6>
        + WAIT_CNT<7> net044 CNT_RST CNT_RST' VDD VSS asynccounter_8
    Xi26 CLK net049 net052 VDD VSS nand2
    Xi19 WAIT_CNT<7> CONF_WAITCYCLES<7> WAITHIGH<7> VDD VSS nand2
    Xi18 WAIT_CNT<6> CONF_WAITCYCLES<6> WAITHIGH<6> VDD VSS nand2
    Xi17 WAIT_CNT<5> CONF_WAITCYCLES<5> WAITHIGH<5> VDD VSS nand2
    Xi10 WAIT_CNT<4> CONF_WAITCYCLES<4> WAITHIGH<4> VDD VSS nand2
    Xi3 WAIT_CNT<3> CONF_WAITCYCLES<3> WAITHIGH<3> VDD VSS nand2
    Xi2 WAIT_CNT<2> CONF_WAITCYCLES<2> WAITHIGH<2> VDD VSS nand2
    Xi1 WAIT_CNT<1> CONF_WAITCYCLES<1> WAITHIGH<1> VDD VSS nand2
    Xi0 WAIT_CNT<0> CONF_WAITCYCLES<0> WAITHIGH<0> VDD VSS nand2
    Xi15 net14 net13 WAIT_RST_RST' VDD VSS nand2
    Xi11 net19 net18 WAIT_RST VDD VSS nand2
    Xi5 WAIT_RST' RST' CNT_RST VDD VSS nand2
    Xi22 net025 net030 net029 VDD VSS nor2
    Xi12 EDGE EDGE' WAIT_RST' VDD VSS nor2
    Xi6 WAIT_RST RST CNT_RST' VDD VSS nor2
    Xi25 ENABLE_E2L net049 net050 RST RST' VDD VSS dff_st_ar_dh
    Xi24 READY WAIT_READY net034 RST RST' VDD VSS dff_st_ar_dh
    Xi8 INT EDGE net18 WAIT_RST_RST WAIT_RST_RST' VDD VSS dff_st_ar_dh
    Xi7 net15 EDGE' net19 WAIT_RST_RST WAIT_RST_RST' VDD VSS dff_st_ar_dh
    Xi23 net029 READY VDD VSS inv
    Xi16 WAIT_RST_RST' WAIT_RST_RST VDD VSS inv
    Xi9 INT net15 VDD VSS inv
    Xi14 WAIT_CNT<4> WAIT_CNT<5> WAIT_CNT<6> WAIT_CNT<7> net13 VDD VSS nor4
    Xi13 WAIT_CNT<0> WAIT_CNT<1> WAIT_CNT<2> WAIT_CNT<3> net14 VDD VSS nor4
    Xi21 WAITHIGH<0> WAITHIGH<1> WAITHIGH<2> WAITHIGH<3> net025 VDD VSS nand4
    Xi20 WAITHIGH<4> WAITHIGH<5> WAITHIGH<6> WAITHIGH<7> net030 VDD VSS nand4
    Xi27 net052 CLK_INT VDD VSS buffer
.ENDS

.SUBCKT tdc_ready_v0 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
                     + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6>
                     + CONF_MAXCYCLES<7> CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2>
                     + CONF_WAITCYCLES<3> CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                     + CONF_WAITCYCLES<7> ENABLE_E2L FF0<0> FF0<1> FF0<2> FF1<0> FF1<1> FF1<2> INT
                     + READY RST RST' VDD VSS
    Xi18 FF0<0> FF0<1> FF0<2> FF1<0> FF1<1> FF1<2> FF_Ready RST RST' VDD VSS ff_ready
    Xi20 CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4>
         + CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> INT net017 RST RST' VDD VSS
         + max_ready
    Xi32 ALARM<0> net19 net027 READY_I VDD VSS nand3
    Xi19 CLK CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
         + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
         + INT RST RST' VDD VSS WAIT_Ready wait_ready
    Xi28 WAIT_Ready net19 VDD VSS inv
    Xi27 FF_Ready ALARM<0> VDD VSS inv
    Xi30 READY_I READY Ready' RST RST' VDD VSS dff_st_ar_dh
    Xi33 net017 Ready' ALARM<1> net027 RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT tdc_and_diff IN0_N IN0_P IN1_N IN1_P OUT_N OUT_P VDD VSS
    Mm3 net18 IN1_P VSS VSS n_mos l=60n w=240.0n m=1
    Mm2 OUT_N IN0_P net18 VSS n_mos l=60n w=240.0n m=1
    Mm1 OUT_P IN0_N VSS VSS n_mos l=60n w=120.0n m=1
    Mm0 OUT_P IN1_N VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 OUT_N OUT_P VDD VDD p_mos l=60n w=120.0n m=1
    Mm4 OUT_P OUT_N VDD VDD p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_buf_diff_np_4lin CONF_N<0> CONF_N<1> CONF_N<2> CONF_N<3> CONF_P<0> CONF_P<1> CONF_P<2>
                             + CONF_P<3> IN_N IN_P OUT_N OUT_P VDD VSS
    Mm51 CONF_N'<3> CONF_N<3> VSS VSS n_mos l=60n w=120.0n m=1
    Mm50 CONF_N'<2> CONF_N<2> VSS VSS n_mos l=60n w=120.0n m=1
    Mm49 CONF_N'<1> CONF_N<1> VSS VSS n_mos l=60n w=120.0n m=1
    Mm48 CONF_N'<0> CONF_N<0> VSS VSS n_mos l=60n w=120.0n m=1
    Mm43 CONF_P'<3> CONF_P<3> VSS VSS n_mos l=60n w=120.0n m=1
    Mm42 CONF_P'<2> CONF_P<2> VSS VSS n_mos l=60n w=120.0n m=1
    Mm41 CONF_P'<1> CONF_P<1> VSS VSS n_mos l=60n w=120.0n m=1
    Mm40 CONF_P'<0> CONF_P<0> VSS VSS n_mos l=60n w=120.0n m=1
    Mm35 OUT_P IN_N VSS VSS n_mos l=60n w=120.0n m=1
    Mm33 OUT_N IN_P VSS VSS n_mos l=60n w=120.0n m=1
    Mm15 net49 CONF_N<3> VSS VSS n_mos l=60n w=120.0n m=1
    Mm14 net52 CONF_N<2> VSS VSS n_mos l=60n w=120.0n m=1
    Mm13 net53 CONF_N<1> VSS VSS n_mos l=60n w=120.0n m=1
    Mm12 net56 CONF_N<0> VSS VSS n_mos l=60n w=120.0n m=1
    Mm11 OUT_P OUT_N net49 VSS n_mos l=60n w=120.0n m=1
    Mm10 OUT_P OUT_N net52 VSS n_mos l=60n w=120.0n m=1
    Mm9 OUT_P OUT_N net53 VSS n_mos l=60n w=120.0n m=1
    Mm8 OUT_P OUT_N net56 VSS n_mos l=60n w=120.0n m=1
    Mm7 net57 CONF_P<3> VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 net60 CONF_P<2> VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 net61 CONF_P<1> VSS VSS n_mos l=60n w=120.0n m=1
    Mm4 net64 CONF_P<0> VSS VSS n_mos l=60n w=120.0n m=1
    Mm3 OUT_N OUT_P net57 VSS n_mos l=60n w=120.0n m=1
    Mm2 OUT_N OUT_P net60 VSS n_mos l=60n w=120.0n m=1
    Mm1 OUT_N OUT_P net61 VSS n_mos l=60n w=120.0n m=1
    Mm0 OUT_N OUT_P net64 VSS n_mos l=60n w=120.0n m=1
    Mm47 CONF_N'<3> CONF_N<3> VDD VDD p_mos l=60n w=120.0n m=1
    Mm46 CONF_N'<2> CONF_N<2> VDD VDD p_mos l=60n w=120.0n m=1
    Mm45 CONF_N'<1> CONF_N<1> VDD VDD p_mos l=60n w=120.0n m=1
    Mm44 CONF_N'<0> CONF_N<0> VDD VDD p_mos l=60n w=120.0n m=1
    Mm39 CONF_P'<3> CONF_P<3> VDD VDD p_mos l=60n w=120.0n m=1
    Mm38 CONF_P'<2> CONF_P<2> VDD VDD p_mos l=60n w=120.0n m=1
    Mm37 CONF_P'<1> CONF_P<1> VDD VDD p_mos l=60n w=120.0n m=1
    Mm36 CONF_P'<0> CONF_P<0> VDD VDD p_mos l=60n w=120.0n m=1
    Mm34 OUT_P IN_N VDD VDD p_mos l=60n w=120.0n m=1
    Mm32 OUT_N IN_P VDD VDD p_mos l=60n w=120.0n m=1
    Mm31 OUT_P OUT_N net50 VDD p_mos l=60n w=120.0n m=1
    Mm30 OUT_P OUT_N net51 VDD p_mos l=60n w=120.0n m=1
    Mm29 OUT_P OUT_N net54 VDD p_mos l=60n w=120.0n m=1
    Mm28 OUT_P OUT_N net55 VDD p_mos l=60n w=120.0n m=1
    Mm27 net50 CONF_P'<3> VDD VDD p_mos l=60n w=120.0n m=1
    Mm26 net51 CONF_P'<2> VDD VDD p_mos l=60n w=120.0n m=1
    Mm25 net54 CONF_P'<1> VDD VDD p_mos l=60n w=120.0n m=1
    Mm24 net55 CONF_P'<0> VDD VDD p_mos l=60n w=120.0n m=1
    Mm23 OUT_N OUT_P net58 VDD p_mos l=60n w=120.0n m=1
    Mm22 OUT_N OUT_P net59 VDD p_mos l=60n w=120.0n m=1
    Mm21 OUT_N OUT_P net62 VDD p_mos l=60n w=120.0n m=1
    Mm20 OUT_N OUT_P net63 VDD p_mos l=60n w=120.0n m=1
    Mm19 net58 CONF_N'<3> VDD VDD p_mos l=60n w=120.0n m=1
    Mm18 net59 CONF_N'<2> VDD VDD p_mos l=60n w=120.0n m=1
    Mm17 net62 CONF_N'<1> VDD VDD p_mos l=60n w=120.0n m=1
    Mm16 net63 CONF_N'<0> VDD VDD p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_inv IN OUT VDD VSS
    Mm0 OUT IN VDD VDD p_mos l=60n w=120.0n m=1
    Mm1 OUT IN VSS VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_inv_wide IN OUT VDD VSS
    Mm0 OUT IN VSS VSS n_mos l=60n w=480.0n m=1
    Mm1 OUT IN VDD VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT tdc_stage_diff_np_4lin_buf CONF_N<0> CONF_N<1> CONF_N<2> CONF_N<3> CONF_P<0> CONF_P<1>
                                   + CONF_P<2> CONF_P<3> IN0_N IN0_P IN1_N IN1_P OUT_BUF_N OUT_BUF_P
                                   + OUT_N OUT_P VDD VSS
    Xi0 IN0_N IN0_P IN1_N IN1_P INT_N INT_P VDD VSS tdc_and_diff
    Xi1 CONF_N<0> CONF_N<1> CONF_N<2> CONF_N<3> CONF_P<0> CONF_P<1> CONF_P<2> CONF_P<3> INT_N INT_P
        + OUT_N_I OUT_P_I VDD VSS tdc_buf_diff_np_4lin
    Xi3 OUT_N OUT_BUF_P VDD VSS tdc_inv
    Xi2 OUT_P OUT_BUF_N VDD VSS tdc_inv
    Xi4 OUT_N_I OUT_P VDD VSS tdc_inv_wide
    Xi5 OUT_P_I OUT_N VDD VSS tdc_inv_wide
.ENDS

.SUBCKT tdc_2stage_diff_np_4lin_buf BUF0_N BUF0_P BUF1_N BUF1_P CONF0_N<0> CONF0_N<1> CONF0_N<2>
                                    + CONF0_N<3> CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3>
                                    + CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_P<0>
                                    + CONF1_P<1> CONF1_P<2> CONF1_P<3> FF0 FF1 IN0_N IN0_P IN1_N
                                    + IN1_P NAND0_IN NAND0_OUT NAND1_IN NAND1_OUT OUT0_N OUT0_P
                                    + OUT1_N OUT1_P RST RST' VDD VSS
    Xi19 OUT_BUF1_N BUF1_N VDD VSS inv_wn
    Xi16 OUT_BUF0_P BUF0_P VDD VSS inv_wn
    Xi17 OUT_BUF0_N BUF0_N VDD VSS inv_wn
    Xi18 OUT_BUF1_P BUF1_P VDD VSS inv_wn
    Xi13 NOR0 NAND0 FF0 Q0' RST RST' VDD VSS dff_st_ar
    Xi12 NOR1 NAND1 FF1 Q1' RST RST' VDD VSS dff_st_ar
    Xi10 Q0' ENABLE0 NAND0_OUT VDD VSS nand2
    Xi11 Q1' ENABLE1 NAND1_OUT VDD VSS nand2
    Xi6 Q1' OUT_BUF0_N NAND1 VDD VSS nand2
    Xi7 Q0' OUT_BUF1_P NAND0 VDD VSS nand2
    Xi9 OUT_BUF0_P NAND0_IN NOR0 VDD VSS nor2
    Xi8 OUT_BUF1_N NAND1_IN NOR1 VDD VSS nor2
    Xi15 NAND0_IN ENABLE0 VDD VSS inv
    Xi14 NAND1_IN ENABLE1 VDD VSS inv
    Xi1 CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3>
        + IN1_N IN1_P NAND1_IN ENABLE1 OUT_BUF1_N OUT_BUF1_P OUT1_N OUT1_P VDD VSS
        + tdc_stage_diff_np_4lin_buf
    Xi0 CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3>
        + IN0_N IN0_P NAND0_IN ENABLE0 OUT_BUF0_N OUT_BUF0_P OUT0_N OUT0_P VDD VSS
        + tdc_stage_diff_np_4lin_buf
.ENDS

.SUBCKT tdc_stage_diff_np_4lin_switched_buf CONF_N<0> CONF_N<1> CONF_N<2> CONF_N<3> CONF_P<0>
                                            + CONF_P<1> CONF_P<2> CONF_P<3> IN0_N IN0_P IN1_N IN1_P
                                            + OUT_BUF_N OUT_BUF_P OUT_N OUT_P VDD VSS
    Xi0 IN0_N IN0_P IN1_N IN1_P INT_N INT_P VDD VSS tdc_and_diff
    Xi1 CONF_N<0> CONF_N<1> CONF_N<2> CONF_N<3> CONF_P<0> CONF_P<1> CONF_P<2> CONF_P<3> INT_P INT_N
        + OUT_N_I OUT_P_I VDD VSS tdc_buf_diff_np_4lin
    Xi3 OUT_N OUT_BUF_P VDD VSS tdc_inv
    Xi2 OUT_P OUT_BUF_N VDD VSS tdc_inv
    Xi4 OUT_N_I OUT_P VDD VSS tdc_inv_wide
    Xi5 OUT_P_I OUT_N VDD VSS tdc_inv_wide
.ENDS

.SUBCKT tdc_2stage_diff_np_4lin_switched_buf BUF0_N BUF0_P BUF1_N BUF1_P CONF0_N<0> CONF0_N<1>
                                             + CONF0_N<2> CONF0_N<3> CONF0_P<0> CONF0_P<1>
                                             + CONF0_P<2> CONF0_P<3> CONF1_N<0> CONF1_N<1>
                                             + CONF1_N<2> CONF1_N<3> CONF1_P<0> CONF1_P<1>
                                             + CONF1_P<2> CONF1_P<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P
                                             + FF0 FF1 IN0_N IN0_P IN1_N IN1_P NAND0_IN NAND0_OUT
                                             + NAND1_IN NAND1_OUT OUT0_N OUT0_P OUT1_N OUT1_P RST
                                             + RST' VDD VSS
    Xi15 NAND1_IN RST' net059 VDD VSS nand2
    Xi14 NAND0_IN RST' net036 VDD VSS nand2
    Xi11 Q1' net059 NAND1_OUT VDD VSS nand2
    Xi10 Q0' net036 NAND0_OUT VDD VSS nand2
    Xi4 Q0' OUT_BUF1_P NAND0 VDD VSS nand2
    Xi5 Q1' OUT_BUF0_N NAND1 VDD VSS nand2
    Xi6 OUT_BUF0_P NAND0_IN NOR0 VDD VSS nor2
    Xi7 OUT_BUF1_N NAND1_IN NOR1 VDD VSS nor2
    Xi8 NOR0 NAND0 FF0 Q0' RST RST' VDD VSS dff_st_ar
    Xi9 NOR1 NAND1 FF1 Q1' RST RST' VDD VSS dff_st_ar
    Xi19 OUT_BUF1_N BUF1_N VDD VSS inv_wn
    Xi18 OUT_BUF1_P BUF1_P VDD VSS inv_wn
    Xi17 OUT_BUF0_N BUF0_N VDD VSS inv_wn
    Xi16 OUT_BUF0_P BUF0_P VDD VSS inv_wn
    Xi1 CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3>
        + IN1_N IN1_P EDGE1_N EDGE1_P OUT_BUF1_N OUT_BUF1_P OUT1_N OUT1_P VDD VSS
        + tdc_stage_diff_np_4lin_switched_buf
    Xi0 CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3>
        + IN0_N IN0_P EDGE0_N EDGE0_P OUT_BUF0_N OUT_BUF0_P OUT0_N OUT0_P VDD VSS
        + tdc_stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT tdc_2e_2b_diff_np_4lin_buf BUF0_N<0> BUF0_N<1> BUF0_N<2> BUF0_P<0> BUF0_P<1> BUF0_P<2>
                                   + BUF1_N<0> BUF1_N<1> BUF1_N<2> BUF1_P<0> BUF1_P<1> BUF1_P<2>
                                   + CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_N<4>
                                   + CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8> CONF0_N<9>
                                   + CONF0_N<10> CONF0_N<11> CONF0_P<0> CONF0_P<1> CONF0_P<2>
                                   + CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7>
                                   + CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<0>
                                   + CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4> CONF1_N<5>
                                   + CONF1_N<6> CONF1_N<7> CONF1_N<8> CONF1_N<9> CONF1_N<10>
                                   + CONF1_N<11> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3>
                                   + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                                   + CONF1_P<9> CONF1_P<10> CONF1_P<11> EDGE0_N EDGE0_P EDGE1_N
                                   + EDGE1_P FF0<0> FF0<1> FF0<2> FF1<0> FF1<1> FF1<2> RST RST' VDD
                                   + VSS
    Xi14 BUF0_N<2> BUF0_P<2> BUF1_N<2> BUF1_P<2> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11>
         + CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<8> CONF1_N<9> CONF1_N<10>
         + CONF1_N<11> CONF1_P<8> CONF1_P<9> CONF1_P<10> CONF1_P<11> FF0<2> FF1<2> INT0_N<1>
         + INT0_P<1> INT1_N<1> INT1_P<1> NAND0<1> NAND0<2> NAND1<1> NAND1<2> INT0_N<2> INT0_P<2>
         + INT1_N<2> INT1_P<2> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi13 BUF0_N<1> BUF0_P<1> BUF1_N<1> BUF1_P<1> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7>
         + CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
         + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> FF0<1> FF1<1> INT0_N<0> INT0_P<0> INT1_N<0>
         + INT1_P<0> NAND0<0> NAND0<1> NAND1<0> NAND1<1> INT0_N<1> INT0_P<1> INT1_N<1> INT1_P<1> RST
         + RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi12 BUF0_N<0> BUF0_P<0> BUF1_N<0> BUF1_P<0> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
         + CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3>
         + CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0> FF1<0>
         + INT1_N<2> INT1_P<2> INT0_N<2> INT0_P<2> NAND1<2> NAND0<0> NAND0<2> NAND1<0> INT0_N<0>
         + INT0_P<0> INT1_N<0> INT1_P<0> RST RST' VDD VSS tdc_2stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT tdc_2b_diff_branch ALARM<0> ALARM<1> BUF1_P<0> CLK CONF0_N<0> CONF0_N<1> CONF0_N<2>
                           + CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8>
                           + CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_P<0> CONF0_P<1> CONF0_P<2>
                           + CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF0_P<8>
                           + CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<0> CONF1_N<1> CONF1_N<2>
                           + CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8>
                           + CONF1_N<9> CONF1_N<10> CONF1_N<11> CONF1_P<0> CONF1_P<1> CONF1_P<2>
                           + CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                           + CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF_DEC<0> CONF_DEC<1> CONF_DEC<2>
                           + CONF_DEC<3> CONF_DEC<4> CONF_DEC<5> CONF_MAXCYCLES<0> CONF_MAXCYCLES<1>
                           + CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5>
                           + CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> CONF_WAITCYCLES<0>
                           + CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
                           + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                           + CONF_WAITCYCLES<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L FF<0>
                           + FF<1> FF<2> FF<3> FF<4> FF<5> RAND_OUT READY RST RST' VDD VSS
    Xi7 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5> FF<0> FF<1> FF<2>
        + FF<3> FF<4> FF<5> RAND_OUT VDD VSS dec_6_conf_0
    Xi2 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
        + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7>
        + CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
        + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
        + FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> BUF0_P<0> READY RST RST' VDD VSS tdc_ready_v0
    Xi1 net025<0> net025<1> net025<2> BUF0_P<0> BUF0_P<1> BUF0_P<2> net024<0> net024<1> net024<2>
        + BUF1_P<0> BUF1_P<1> BUF1_P<2> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_N<4>
        + CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_P<0>
        + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF0_P<8>
        + CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4>
        + CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8> CONF1_N<9> CONF1_N<10> CONF1_N<11> CONF1_P<0>
        + CONF1_P<1> CONF1_P<2> CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
        + CONF1_P<9> CONF1_P<10> CONF1_P<11> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF<0> FF<1> FF<2> FF<3>
        + FF<4> FF<5> RST RST' VDD VSS tdc_2e_2b_diff_np_4lin_buf
.ENDS

.SUBCKT tdc_2e_3b_diff_np_4lin_buf BUF0_N<0> BUF0_N<1> BUF0_N<2> BUF0_N<3> BUF0_P<0> BUF0_P<1>
                                   + BUF0_P<2> BUF0_P<3> BUF1_N<0> BUF1_N<1> BUF1_N<2> BUF1_N<3>
                                   + BUF1_P<0> BUF1_P<1> BUF1_P<2> BUF1_P<3> CONF0_N<0> CONF0_N<1>
                                   + CONF0_N<2> CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6>
                                   + CONF0_N<7> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11>
                                   + CONF0_N<12> CONF0_N<13> CONF0_N<14> CONF0_N<15> CONF0_P<0>
                                   + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5>
                                   + CONF0_P<6> CONF0_P<7> CONF0_P<8> CONF0_P<9> CONF0_P<10>
                                   + CONF0_P<11> CONF0_P<12> CONF0_P<13> CONF0_P<14> CONF0_P<15>
                                   + CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4>
                                   + CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8> CONF1_N<9>
                                   + CONF1_N<10> CONF1_N<11> CONF1_N<12> CONF1_N<13> CONF1_N<14>
                                   + CONF1_N<15> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3>
                                   + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                                   + CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12> CONF1_P<13>
                                   + CONF1_P<14> CONF1_P<15> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0>
                                   + FF0<1> FF0<2> FF0<3> FF1<0> FF1<1> FF1<2> FF1<3> RST RST' VDD
                                   + VSS
    Xi13 BUF0_N<1> BUF0_P<1> BUF1_N<1> BUF1_P<1> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7>
         + CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
         + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> FF0<1> FF1<1> INT0_N<0> INT0_P<0> INT1_N<0>
         + INT1_P<0> NAND0<0> NAND0<1> NAND1<0> NAND1<1> INT0_N<1> INT0_P<1> INT1_N<1> INT1_P<1> RST
         + RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi14 BUF0_N<2> BUF0_P<2> BUF1_N<2> BUF1_P<2> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11>
         + CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<8> CONF1_N<9> CONF1_N<10>
         + CONF1_N<11> CONF1_P<8> CONF1_P<9> CONF1_P<10> CONF1_P<11> FF0<2> FF1<2> INT0_N<1>
         + INT0_P<1> INT1_N<1> INT1_P<1> NAND0<1> NAND0<2> NAND1<1> NAND1<2> INT0_N<2> INT0_P<2>
         + INT1_N<2> INT1_P<2> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi17 BUF0_N<3> BUF0_P<3> BUF1_N<3> BUF1_P<3> CONF0_N<12> CONF0_N<13> CONF0_N<14> CONF0_N<15>
         + CONF0_P<12> CONF0_P<13> CONF0_P<14> CONF0_P<15> CONF1_N<12> CONF1_N<13> CONF1_N<14>
         + CONF1_N<15> CONF1_P<12> CONF1_P<13> CONF1_P<14> CONF1_P<15> FF0<3> FF1<3> INT0_N<2>
         + INT0_P<2> INT1_N<2> INT1_P<2> NAND0<2> NAND0<3> NAND1<2> NAND1<3> INT0_N<3> INT0_P<3>
         + INT1_N<3> INT1_P<3> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi12 BUF0_N<0> BUF0_P<0> BUF1_N<0> BUF1_P<0> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
         + CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3>
         + CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0> FF1<0>
         + INT1_N<3> INT1_P<3> INT0_N<3> INT0_P<3> NAND1<3> NAND0<0> NAND0<3> NAND1<0> INT0_N<0>
         + INT0_P<0> INT1_N<0> INT1_P<0> RST RST' VDD VSS tdc_2stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT ff_ready_4 FF0<0> FF0<1> FF0<2> FF0<3> FF1<0> FF1<1> FF1<2> FF1<3> FF_READY RST RST' VDD VSS
    Xi2 FF_NOR0 FF_NOR1 FF_NAND VDD VSS nand2
    Xi3 FF_NAND FF_READY net18 RST RST' VDD VSS dff_st_ar_dh
    Xi0 FF0<0> FF0<1> FF0<2> FF0<3> FF_NOR0 VDD VSS nor4
    Xi1 FF1<0> FF1<1> FF1<2> FF1<3> FF_NOR1 VDD VSS nor4
.ENDS

.SUBCKT tdc_ready_4 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
                    + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6>
                    + CONF_MAXCYCLES<7> CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2>
                    + CONF_WAITCYCLES<3> CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                    + CONF_WAITCYCLES<7> ENABLE_E2L FF0<0> FF0<1> FF0<2> FF0<3> FF1<0> FF1<1> FF1<2>
                    + FF1<3> INT READY RST RST' VDD VSS
    Xi20 CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4>
         + CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> INT net017 RST RST' VDD VSS
         + max_ready
    Xi32 ALARM<0> net19 net027 READY_I VDD VSS nand3
    Xi19 CLK CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
         + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
         + INT RST RST' VDD VSS WAIT_Ready wait_ready
    Xi28 WAIT_Ready net19 VDD VSS inv
    Xi27 FF_Ready ALARM<0> VDD VSS inv
    Xi30 READY_I READY Ready' RST RST' VDD VSS dff_st_ar_dh
    Xi33 net017 Ready' ALARM<1> net027 RST RST' VDD VSS dff_st_ar
    Xi18 FF0<0> FF0<1> FF0<2> FF0<3> FF1<0> FF1<1> FF1<2> FF1<3> FF_Ready RST RST' VDD VSS
         + ff_ready_4
.ENDS

.SUBCKT dec_8_conf_0 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5>
                     + CONF_DEC<6> CONF_DEC<7> FF_IN<0> FF_IN<1> FF_IN<2> FF_IN<3> FF_IN<4> FF_IN<5>
                     + FF_IN<6> FF_IN<7> RAND_OUT VDD VSS
    Xi28 CONF_DEC<7> FF_IN<7> FF_IN<6> STAGE<7> VDD VSS dec_stage
    Xi27 CONF_DEC<6> FF_IN<6> FF_IN<5> STAGE<6> VDD VSS dec_stage
    Xi23 CONF_DEC<5> FF_IN<5> FF_IN<4> STAGE<5> VDD VSS dec_stage
    Xi22 CONF_DEC<4> FF_IN<4> FF_IN<3> STAGE<4> VDD VSS dec_stage
    Xi21 CONF_DEC<3> FF_IN<3> FF_IN<2> STAGE<3> VDD VSS dec_stage
    Xi20 CONF_DEC<2> FF_IN<2> FF_IN<1> STAGE<2> VDD VSS dec_stage
    Xi19 CONF_DEC<1> FF_IN<1> FF_IN<0> STAGE<1> VDD VSS dec_stage
    Xi18 CONF_DEC<0> FF_IN<0> FF_IN<7> STAGE<0> VDD VSS dec_stage
    Xi26 net026 net023 RAND_OUT VDD VSS nor2
    Xi25 STAGE<4> STAGE<5> STAGE<6> STAGE<7> net023 VDD VSS nand4
    Xi24 STAGE<0> STAGE<1> STAGE<2> STAGE<3> net026 VDD VSS nand4
.ENDS

.SUBCKT tdc_3b_diff_branch ALARM<0> ALARM<1> BUF1_P<0> CLK CONF0_N<0> CONF0_N<1> CONF0_N<2>
                           + CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8>
                           + CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_N<12> CONF0_N<13> CONF0_N<14>
                           + CONF0_N<15> CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4>
                           + CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF0_P<8> CONF0_P<9> CONF0_P<10>
                           + CONF0_P<11> CONF0_P<12> CONF0_P<13> CONF0_P<14> CONF0_P<15> CONF1_N<0>
                           + CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6>
                           + CONF1_N<7> CONF1_N<8> CONF1_N<9> CONF1_N<10> CONF1_N<11> CONF1_N<12>
                           + CONF1_N<13> CONF1_N<14> CONF1_N<15> CONF1_P<0> CONF1_P<1> CONF1_P<2>
                           + CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                           + CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12> CONF1_P<13> CONF1_P<14>
                           + CONF1_P<15> CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4>
                           + CONF_DEC<5> CONF_DEC<6> CONF_DEC<7> CONF_MAXCYCLES<0> CONF_MAXCYCLES<1>
                           + CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5>
                           + CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> CONF_WAITCYCLES<0>
                           + CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
                           + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                           + CONF_WAITCYCLES<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L FF<0>
                           + FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> RAND_OUT READY RST RST' VDD
                           + VSS
    Xi1 net31<0> net31<1> net31<2> net31<3> BUF0_P<0> BUF0_P<1> BUF0_P<2> BUF0_P<3> net30<0>
        + net30<1> net30<2> net30<3> BUF1_P<0> BUF1_P<1> BUF1_P<2> BUF1_P<3> CONF0_N<0> CONF0_N<1>
        + CONF0_N<2> CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8> CONF0_N<9>
        + CONF0_N<10> CONF0_N<11> CONF0_N<12> CONF0_N<13> CONF0_N<14> CONF0_N<15> CONF0_P<0>
        + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF0_P<8>
        + CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF0_P<12> CONF0_P<13> CONF0_P<14> CONF0_P<15>
        + CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
        + CONF1_N<8> CONF1_N<9> CONF1_N<10> CONF1_N<11> CONF1_N<12> CONF1_N<13> CONF1_N<14>
        + CONF1_N<15> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6>
        + CONF1_P<7> CONF1_P<8> CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12> CONF1_P<13>
        + CONF1_P<14> CONF1_P<15> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF<0> FF<1> FF<2> FF<3> FF<4>
        + FF<5> FF<6> FF<7> RST RST' VDD VSS tdc_2e_3b_diff_np_4lin_buf
    Xi2 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
        + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7>
        + CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
        + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
        + FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> BUF0_P<0> READY RST RST' VDD VSS
        + tdc_ready_4
    Xi7 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5> CONF_DEC<6>
        + CONF_DEC<7> FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> RAND_OUT VDD VSS dec_8_conf_0
.ENDS

.SUBCKT dff_st_ar_buf CLK D Q Q' RST RST' VDD VSS
    Xi0 CLK D net17 net18 RST RST' VDD VSS dff_st_ar
    Xi2 net17 Q' VDD VSS inv
    Xi1 net18 Q VDD VSS inv
.ENDS

.SUBCKT edge2level_3e EDGE ENABLE OUT0 OUT1 OUT2 RST RST' VDD VSS
    Xi5 EDGE OUT1 OUT2 net17 RST RST' VDD VSS dff_st_ar_buf
    Xi4 EDGE OUT0 OUT1 net18 RST RST' VDD VSS dff_st_ar_buf
    Xi3 EDGE ENABLE OUT0 net19 RST RST' VDD VSS dff_st_ar_buf
.ENDS

.SUBCKT mero_nand2 IN0 IN1 OUT VDD VSS
    Mm1 OUT IN1 VDD VDD p_mos l=60n w=120.0n m=1
    Mm0 OUT IN0 VDD VDD p_mos l=60n w=120.0n m=1
    Mm3 net7 IN1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm2 OUT IN0 net7 VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT mero_buf IN OUT VDD VSS
    Mm1 OUT net1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm0 net1 IN VSS VSS n_mos l=60n w=120.0n m=1
    Mm3 OUT net1 VDD VDD p_mos l=60n w=120.0n m=1
    Mm2 net1 IN VDD VDD p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT mero_3e_1b ENABLE OUT0 OUT1 OUT2 VDD VSS
    Xi2 OUT1 ENABLE net5 VDD VSS mero_nand2
    Xi1 OUT0 ENABLE net6 VDD VSS mero_nand2
    Xi0 OUT2 ENABLE net7 VDD VSS mero_nand2
    Xi5 net5 OUT2 VDD VSS mero_buf
    Xi4 net6 OUT1 VDD VSS mero_buf
    Xi3 net7 OUT0 VDD VSS mero_buf
.ENDS

.SUBCKT dc_3e_1b_noconfig ENABLE_E2L ENABLE_MERO INT0 INT1 INT2 OUT0 OUT1 OUT2 RST RST' VDD VSS
    Xi11 MERO_OUT2 INT2 VDD VSS buffer
    Xi9 MERO_OUT0 INT0 VDD VSS buffer
    Xi10 MERO_OUT1 INT1 VDD VSS buffer
    Xi1 INT1 ENABLE_E2L OUT0 OUT1 OUT2 RST RST' VDD VSS edge2level_3e
    Xi5 ENABLE_INT MERO_OUT0 MERO_OUT1 MERO_OUT2 VDD VSS mero_3e_1b
    Xi12 OUT2 net10 ENABLE_INT VDD VSS nor2
    Xi13 ENABLE_MERO net10 VDD VSS inv
.ENDS

.SUBCKT mero_3e_4b ENABLE OUT0 OUT1 OUT2 VDD VSS
    Xi2 OUT1 ENABLE INT2<0> VDD VSS mero_nand2
    Xi1 OUT0 ENABLE INT1<0> VDD VSS mero_nand2
    Xi0 OUT2 ENABLE INT0<0> VDD VSS mero_nand2
    Xi14 INT2<3> OUT2 VDD VSS mero_buf
    Xi13 INT1<3> OUT1 VDD VSS mero_buf
    Xi12 INT0<3> OUT0 VDD VSS mero_buf
    Xi11 INT2<2> INT2<3> VDD VSS mero_buf
    Xi10 INT1<2> INT1<3> VDD VSS mero_buf
    Xi9 INT0<2> INT0<3> VDD VSS mero_buf
    Xi8 INT2<1> INT2<2> VDD VSS mero_buf
    Xi7 INT2<0> INT2<1> VDD VSS mero_buf
    Xi6 INT1<1> INT1<2> VDD VSS mero_buf
    Xi5 INT1<0> INT1<1> VDD VSS mero_buf
    Xi4 INT0<1> INT0<2> VDD VSS mero_buf
    Xi3 INT0<0> INT0<1> VDD VSS mero_buf
.ENDS

.SUBCKT dc_3e_4b_noconfig ENABLE_E2L ENABLE_MERO INT0 INT1 INT2 OUT0 OUT1 OUT2 RST RST' VDD VSS
    Xi11 MERO_OUT2 INT2 VDD VSS buffer
    Xi9 MERO_OUT0 INT0 VDD VSS buffer
    Xi10 MERO_OUT1 INT1 VDD VSS buffer
    Xi1 INT1 ENABLE_E2L OUT0 OUT1 OUT2 RST RST' VDD VSS edge2level_3e
    Xi5 ENABLE_INT MERO_OUT0 MERO_OUT1 MERO_OUT2 VDD VSS mero_3e_4b
    Xi12 OUT2 net013 ENABLE_INT VDD VSS nor2
    Xi13 ENABLE_MERO net013 VDD VSS inv
.ENDS

.SUBCKT mero_3e_3b ENABLE OUT0 OUT1 OUT2 VDD VSS
    Xi2 OUT1 ENABLE INT2<0> VDD VSS mero_nand2
    Xi1 OUT0 ENABLE INT1<0> VDD VSS mero_nand2
    Xi0 OUT2 ENABLE INT0<0> VDD VSS mero_nand2
    Xi14 INT2<2> OUT2 VDD VSS mero_buf
    Xi13 INT1<2> OUT1 VDD VSS mero_buf
    Xi12 INT0<2> OUT0 VDD VSS mero_buf
    Xi8 INT2<1> INT2<2> VDD VSS mero_buf
    Xi7 INT2<0> INT2<1> VDD VSS mero_buf
    Xi6 INT1<1> INT1<2> VDD VSS mero_buf
    Xi5 INT1<0> INT1<1> VDD VSS mero_buf
    Xi4 INT0<1> INT0<2> VDD VSS mero_buf
    Xi3 INT0<0> INT0<1> VDD VSS mero_buf
.ENDS

.SUBCKT dc_3e_3b_noconfig ENABLE_E2L ENABLE_MERO INT0 INT1 INT2 OUT0 OUT1 OUT2 RST RST' VDD VSS
    Xi11 MERO_OUT2 INT2 VDD VSS buffer
    Xi9 MERO_OUT0 INT0 VDD VSS buffer
    Xi10 MERO_OUT1 INT1 VDD VSS buffer
    Xi1 INT1 ENABLE_E2L OUT0 OUT1 OUT2 RST RST' VDD VSS edge2level_3e
    Xi12 OUT2 net014 ENABLE_INT VDD VSS nor2
    Xi5 ENABLE_INT MERO_OUT0 MERO_OUT1 MERO_OUT2 VDD VSS mero_3e_3b
    Xi13 ENABLE_MERO net014 VDD VSS inv
.ENDS

.SUBCKT singleended2diff IN OUT_N OUT_P VDD VSS
    Mm2 OUT_N IN VDD VDD p_mos l=60n w=480.0n m=4
    Mm3 OUT_P OUT_N VDD VDD p_mos l=60n w=480.0n m=4
    Mm1 OUT_P OUT_N VSS VSS n_mos l=60n w=480.0n m=4
    Mm0 OUT_N IN VSS VSS n_mos l=60n w=480.0n m=4
.ENDS

.SUBCKT mux4 IN<0> IN<1> IN<2> IN<3> OUT SEL<0> SEL<1> VDD VSS
    Xi2 net8 net7 OUT SEL<1> VDD VSS mux2
    Xi1 IN<2> IN<3> net7 SEL<0> VDD VSS mux2
    Xi0 IN<0> IN<1> net8 SEL<0> VDD VSS mux2
.ENDS

.SUBCKT dec4_inverted OUT<0> OUT<1> OUT<2> OUT<3> SEL<0> SEL<1> VDD VSS
    Xi1 SEL<1> SEL'<1> VDD VSS inv
    Xi0 SEL<0> SEL'<0> VDD VSS inv
    Xi6 SEL<0> SEL<1> OUT<3> VDD VSS nand2
    Xi5 SEL'<0> SEL<1> OUT<2> VDD VSS nand2
    Xi4 SEL<0> SEL'<1> OUT<1> VDD VSS nand2
    Xi3 SEL'<0> SEL'<1> OUT<0> VDD VSS nand2
.ENDS

.SUBCKT mero_3e_2b ENABLE OUT0 OUT1 OUT2 VDD VSS
    Xi2 OUT1 ENABLE INT2<0> VDD VSS mero_nand2
    Xi1 OUT0 ENABLE INT1<0> VDD VSS mero_nand2
    Xi0 OUT2 ENABLE INT0<0> VDD VSS mero_nand2
    Xi8 INT2<1> OUT2 VDD VSS mero_buf
    Xi7 INT2<0> INT2<1> VDD VSS mero_buf
    Xi6 INT1<1> OUT1 VDD VSS mero_buf
    Xi5 INT1<0> INT1<1> VDD VSS mero_buf
    Xi4 INT0<1> OUT0 VDD VSS mero_buf
    Xi3 INT0<0> INT0<1> VDD VSS mero_buf
.ENDS

.SUBCKT dc_3e_2b_noconfig ENABLE_E2L ENABLE_MERO INT0 INT1 INT2 OUT0 OUT1 OUT2 RST RST' VDD VSS
    Xi5 ENABLE_INT MERO_OUT0 MERO_OUT1 MERO_OUT2 VDD VSS mero_3e_2b
    Xi1 INT1 ENABLE_E2L OUT0 OUT1 OUT2 RST RST' VDD VSS edge2level_3e
    Xi12 OUT2 net014 ENABLE_INT VDD VSS nor2
    Xi9 MERO_OUT0 INT0 VDD VSS buffer
    Xi11 MERO_OUT2 INT2 VDD VSS buffer
    Xi10 MERO_OUT1 INT1 VDD VSS buffer
    Xi13 ENABLE_MERO net014 VDD VSS inv
.ENDS

.SUBCKT xor2 IN0 IN1 OUT VDD VSS
    Mm3 OUT IN0' net20 VDD p_mos l=60n w=240.0n m=1
    Mm2 net20 IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN0 net21 VDD p_mos l=60n w=240.0n m=1
    Mm0 net21 IN1' VDD VDD p_mos l=60n w=240.0n m=1
    Mm7 net19 IN1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 net18 IN1' VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 OUT IN0' net18 VSS n_mos l=60n w=120.0n m=1
    Mm4 OUT IN0 net19 VSS n_mos l=60n w=120.0n m=1
    Xi1 IN1 IN1' VDD VSS inv
    Xi0 IN0 IN0' VDD VSS inv
.ENDS

.SUBCKT mero_collapse_3e_v2 ALARM ENABLE_E2L INT0 INT1 INT2 RST RST' VDD VSS
    Xi2 INT2 INT1 XOR2 VDD VSS xor2
    Xi1 INT0 INT2 XOR1 VDD VSS xor2
    Xi0 INT1 INT0 XOR0 VDD VSS xor2
    Xi7 NOR OR VDD VSS inv
    Xi4 XOR0 XOR1 XOR2 NOR VDD VSS nor3
    Xi6 ENABLE_E2L OR ALARM net016 RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT vdd_gate_1ma ENABLE' VDD_IN VDD_OUT VSS
    Mm0 VDD_OUT ENABLE' VDD_IN VDD_IN pch_lvt l=60n w=4u m=40
    Mm1 VDD_OUT ENABLE' VSS VSS nch_lvt l=60n w=4u m=40
.ENDS

.SUBCKT dc_collection ALARM_DC CONF_SELDC<0> CONF_SELDC<1> DCEDGE0<1> DCEDGE0<2> DCEDGE0<3>
                      + DCEDGE1<1> DCEDGE1<2> DCEDGE1<3> DCEDGE2<1> DCEDGE2<2> DCEDGE2<3> EDGE0_N
                      + EDGE0_P EDGE1_N EDGE1_P EDGE2_N EDGE2_P ENABLE_E2L ENABLE_MERO MERO_INT<0>
                      + MERO_INT<1> MERO_INT<2> RST RST' SEL_DCEDGE<0> SEL_DCEDGE<1> VDD_CORE VDD_DC
                      + VSS
    Xi29 ENABLE_E2L ENABLE_MERO MERO_INT0<0> MERO_INT1<0> MERO_INT2<0> MERO_EDGE0<0> MERO_EDGE1<0>
         + MERO_EDGE2<0> RST RST' VDD_DC_INT<0> VSS dc_3e_1b_noconfig
    Xi27 ENABLE_E2L ENABLE_MERO MERO_INT0<3> MERO_INT1<3> MERO_INT2<3> MERO_EDGE0<3> MERO_EDGE1<3>
         + MERO_EDGE2<3> RST RST' VDD_DC_INT<3> VSS dc_3e_4b_noconfig
    Xi0 ENABLE_E2L ENABLE_MERO MERO_INT0<2> MERO_INT1<2> MERO_INT2<2> MERO_EDGE0<2> MERO_EDGE1<2>
        + MERO_EDGE2<2> RST RST' VDD_DC_INT<2> VSS dc_3e_3b_noconfig
    Xi9 SEDGE0 EDGE0_N EDGE0_P VDD_DC VSS singleended2diff
    Xi11 SEDGE1 EDGE1_N EDGE1_P VDD_DC VSS singleended2diff
    Xi10 SEDGE2 EDGE2_N EDGE2_P VDD_DC VSS singleended2diff
    Xi21 MERO_EDGE0<0> MERO_EDGE0<1> MERO_EDGE0<2> MERO_EDGE0<3> DCEDGE0<0> CONF_SELDC<0>
         + CONF_SELDC<1> VDD_CORE VSS mux4
    Xi19 MERO_INT0<0> MERO_INT0<1> MERO_INT0<2> MERO_INT0<3> MERO_INT<0> CONF_SELDC<0> CONF_SELDC<1>
         + VDD_CORE VSS mux4
    Xi14 DCEDGE0<0> DCEDGE0<1> DCEDGE0<2> DCEDGE0<3> SEDGE0 SEL_DCEDGE<0> SEL_DCEDGE<1> VDD_CORE VSS
         + mux4
    Xi22 MERO_EDGE1<0> MERO_EDGE1<1> MERO_EDGE1<2> MERO_EDGE1<3> DCEDGE1<0> CONF_SELDC<0>
         + CONF_SELDC<1> VDD_CORE VSS mux4
    Xi18 MERO_INT1<0> MERO_INT1<1> MERO_INT1<2> MERO_INT1<3> MERO_INT<1> CONF_SELDC<0> CONF_SELDC<1>
         + VDD_CORE VSS mux4
    Xi15 DCEDGE1<0> DCEDGE1<1> DCEDGE1<2> DCEDGE1<3> SEDGE1 SEL_DCEDGE<0> SEL_DCEDGE<1> VDD_CORE VSS
         + mux4
    Xi20 MERO_EDGE2<0> MERO_EDGE2<1> MERO_EDGE2<2> MERO_EDGE2<3> DCEDGE2<0> CONF_SELDC<0>
         + CONF_SELDC<1> VDD_CORE VSS mux4
    Xi17 MERO_INT2<0> MERO_INT2<1> MERO_INT2<2> MERO_INT2<3> MERO_INT<2> CONF_SELDC<0> CONF_SELDC<1>
         + VDD_CORE VSS mux4
    Xi16 DCEDGE2<0> DCEDGE2<1> DCEDGE2<2> DCEDGE2<3> SEDGE2 SEL_DCEDGE<0> SEL_DCEDGE<1> VDD_CORE VSS
         + mux4
    Xi30 SELDC_DEC<0> SELDC_DEC<1> SELDC_DEC<2> SELDC_DEC<3> CONF_SELDC<0> CONF_SELDC<1> VDD_CORE
         + VSS dec4_inverted
    Xi24 ENABLE_E2L ENABLE_MERO MERO_INT0<1> MERO_INT1<1> MERO_INT2<1> MERO_EDGE0<1> MERO_EDGE1<1>
         + MERO_EDGE2<1> RST RST' VDD_DC_INT<1> VSS dc_3e_2b_noconfig
    Xi3 ALARM_DC ENABLE_E2L MERO_INT<0> MERO_INT<1> MERO_INT<2> RST RST' VDD_DC VSS
        + mero_collapse_3e_v2
    Xi28 SELDC_DEC<0> VDD_DC VDD_DC_INT<0> VSS vdd_gate_1ma
    Xi26 SELDC_DEC<3> VDD_DC VDD_DC_INT<3> VSS vdd_gate_1ma
    Xi25 SELDC_DEC<1> VDD_DC VDD_DC_INT<1> VSS vdd_gate_1ma
    Xi23 SELDC_DEC<2> VDD_DC VDD_DC_INT<2> VSS vdd_gate_1ma
.ENDS

.SUBCKT dec_10_conf_0 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5>
                      + CONF_DEC<6> CONF_DEC<7> CONF_DEC<8> CONF_DEC<9> FF_IN<0> FF_IN<1> FF_IN<2>
                      + FF_IN<3> FF_IN<4> FF_IN<5> FF_IN<6> FF_IN<7> FF_IN<8> FF_IN<9> RAND_OUT VDD
                      + VSS
    Xi30 CONF_DEC<9> FF_IN<9> FF_IN<8> STAGE<9> VDD VSS dec_stage
    Xi28 CONF_DEC<7> FF_IN<7> FF_IN<6> STAGE<7> VDD VSS dec_stage
    Xi27 CONF_DEC<6> FF_IN<6> FF_IN<5> STAGE<6> VDD VSS dec_stage
    Xi23 CONF_DEC<5> FF_IN<5> FF_IN<4> STAGE<5> VDD VSS dec_stage
    Xi22 CONF_DEC<4> FF_IN<4> FF_IN<3> STAGE<4> VDD VSS dec_stage
    Xi21 CONF_DEC<3> FF_IN<3> FF_IN<2> STAGE<3> VDD VSS dec_stage
    Xi20 CONF_DEC<2> FF_IN<2> FF_IN<1> STAGE<2> VDD VSS dec_stage
    Xi19 CONF_DEC<1> FF_IN<1> FF_IN<0> STAGE<1> VDD VSS dec_stage
    Xi18 CONF_DEC<0> FF_IN<0> FF_IN<9> STAGE<0> VDD VSS dec_stage
    Xi29 CONF_DEC<8> FF_IN<8> FF_IN<7> STAGE<8> VDD VSS dec_stage
    Xi31 STAGE<8> STAGE<9> net038 VDD VSS nand2
    Xi25 STAGE<4> STAGE<5> STAGE<6> STAGE<7> net023 VDD VSS nand4
    Xi24 STAGE<0> STAGE<1> STAGE<2> STAGE<3> net026 VDD VSS nand4
    Xi26 net026 net023 net038 RAND_OUT VDD VSS nor3
.ENDS

.SUBCKT tdc_2e_4b_diff_np_4lin_buf BUF0_N<0> BUF0_N<1> BUF0_N<2> BUF0_N<3> BUF0_N<4> BUF0_P<0>
                                   + BUF0_P<1> BUF0_P<2> BUF0_P<3> BUF0_P<4> BUF1_N<0> BUF1_N<1>
                                   + BUF1_N<2> BUF1_N<3> BUF1_N<4> BUF1_P<0> BUF1_P<1> BUF1_P<2>
                                   + BUF1_P<3> BUF1_P<4> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
                                   + CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8>
                                   + CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_N<12> CONF0_N<13>
                                   + CONF0_N<14> CONF0_N<15> CONF0_N<16> CONF0_N<17> CONF0_N<18>
                                   + CONF0_N<19> CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3>
                                   + CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF0_P<8>
                                   + CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF0_P<12> CONF0_P<13>
                                   + CONF0_P<14> CONF0_P<15> CONF0_P<16> CONF0_P<17> CONF0_P<18>
                                   + CONF0_P<19> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3>
                                   + CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8>
                                   + CONF1_N<9> CONF1_N<10> CONF1_N<11> CONF1_N<12> CONF1_N<13>
                                   + CONF1_N<14> CONF1_N<15> CONF1_N<16> CONF1_N<17> CONF1_N<18>
                                   + CONF1_N<19> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3>
                                   + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                                   + CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12> CONF1_P<13>
                                   + CONF1_P<14> CONF1_P<15> CONF1_P<16> CONF1_P<17> CONF1_P<18>
                                   + CONF1_P<19> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0> FF0<1>
                                   + FF0<2> FF0<3> FF0<4> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> RST
                                   + RST' VDD VSS
    Xi21 BUF0_N<2> BUF0_P<2> BUF1_N<2> BUF1_P<2> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11>
         + CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF1_N<8> CONF1_N<9> CONF1_N<10>
         + CONF1_N<11> CONF1_P<8> CONF1_P<9> CONF1_P<10> CONF1_P<11> FF0<2> FF1<2> INT0_N<1>
         + INT0_P<1> INT1_N<1> INT1_P<1> NAND0<1> NAND0<2> NAND1<1> NAND1<2> INT0_N<2> INT0_P<2>
         + INT1_N<2> INT1_P<2> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi20 BUF0_N<1> BUF0_P<1> BUF1_N<1> BUF1_P<1> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7>
         + CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
         + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> FF0<1> FF1<1> INT0_N<0> INT0_P<0> INT1_N<0>
         + INT1_P<0> NAND0<0> NAND0<1> NAND1<0> NAND1<1> INT0_N<1> INT0_P<1> INT1_N<1> INT1_P<1> RST
         + RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi19 BUF0_N<4> BUF0_P<4> BUF1_N<4> BUF1_P<4> CONF0_N<16> CONF0_N<17> CONF0_N<18> CONF0_N<19>
         + CONF0_P<16> CONF0_P<17> CONF0_P<18> CONF0_P<19> CONF1_N<16> CONF1_N<17> CONF1_N<18>
         + CONF1_N<19> CONF1_P<16> CONF1_P<17> CONF1_P<18> CONF1_P<19> FF0<4> FF1<4> INT0_N<3>
         + INT0_P<3> INT1_N<3> INT1_P<3> NAND0<3> NAND0<4> NAND1<3> NAND1<4> INT0_N<4> INT0_P<4>
         + INT1_N<4> INT1_P<4> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi18 BUF0_N<3> BUF0_P<3> BUF1_N<3> BUF1_P<3> CONF0_N<12> CONF0_N<13> CONF0_N<14> CONF0_N<15>
         + CONF0_P<12> CONF0_P<13> CONF0_P<14> CONF0_P<15> CONF1_N<12> CONF1_N<13> CONF1_N<14>
         + CONF1_N<15> CONF1_P<12> CONF1_P<13> CONF1_P<14> CONF1_P<15> FF0<3> FF1<3> INT0_N<2>
         + INT0_P<2> INT1_N<2> INT1_P<2> NAND0<2> NAND0<3> NAND1<2> NAND1<3> INT0_N<3> INT0_P<3>
         + INT1_N<3> INT1_P<3> RST RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi22 BUF0_N<0> BUF0_P<0> BUF1_N<0> BUF1_P<0> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
         + CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3>
         + CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0> FF1<0>
         + INT1_N<4> INT1_P<4> INT0_N<4> INT0_P<4> NAND1<4> NAND0<0> NAND0<4> NAND1<0> INT0_N<0>
         + INT0_P<0> INT1_N<0> INT1_P<0> RST RST' VDD VSS tdc_2stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT nor5 IN0 IN1 IN2 IN3 IN4 OUT VDD VSS
    Mm8 OUT IN0 net011 VDD p_mos l=60n w=480.0n m=1
    Mm3 net011 IN1 net7 VDD p_mos l=60n w=480.0n m=1
    Mm2 net7 IN2 net6 VDD p_mos l=60n w=480.0n m=1
    Mm1 net6 IN3 net5 VDD p_mos l=60n w=480.0n m=1
    Mm0 net5 IN4 VDD VDD p_mos l=60n w=480.0n m=1
    Mm9 OUT IN0 VSS VSS n_mos l=60n w=120.0n m=1
    Mm7 OUT IN4 VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 OUT IN3 VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 OUT IN1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm4 OUT IN2 VSS VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT ff_ready_6 FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF_READY
                   + RST RST' VDD VSS
    Xi0 FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF_NOR0 VDD VSS nor5
    Xi1 FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF_NOR1 VDD VSS nor5
    Xi2 FF_NOR0 FF_NOR1 FF_NAND VDD VSS nand2
    Xi3 FF_NAND FF_READY net18 RST RST' VDD VSS dff_st_ar_dh
.ENDS

.SUBCKT tdc_ready_6 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
                    + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6>
                    + CONF_MAXCYCLES<7> CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2>
                    + CONF_WAITCYCLES<3> CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                    + CONF_WAITCYCLES<7> ENABLE_E2L FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF1<0> FF1<1>
                    + FF1<2> FF1<3> FF1<4> INT READY RST RST' VDD VSS
    Xi18 FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF_Ready RST RST' VDD
         + VSS ff_ready_6
    Xi20 CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4>
         + CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> INT net017 RST RST' VDD VSS
         + max_ready
    Xi32 ALARM<0> net19 net027 READY_I VDD VSS nand3
    Xi19 CLK CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
         + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
         + INT RST RST' VDD VSS WAIT_Ready wait_ready
    Xi28 WAIT_Ready net19 VDD VSS inv
    Xi27 FF_Ready ALARM<0> VDD VSS inv
    Xi30 READY_I READY Ready' RST RST' VDD VSS dff_st_ar_dh
    Xi33 net017 Ready' ALARM<1> net027 RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT tdc_4b_diff_branch ALARM<0> ALARM<1> BUF1_P<0> CLK CONF0_N<0> CONF0_N<1> CONF0_N<2>
                           + CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_N<8>
                           + CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_N<12> CONF0_N<13> CONF0_N<14>
                           + CONF0_N<15> CONF0_N<16> CONF0_N<17> CONF0_N<18> CONF0_N<19> CONF0_P<0>
                           + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6>
                           + CONF0_P<7> CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF0_P<12>
                           + CONF0_P<13> CONF0_P<14> CONF0_P<15> CONF0_P<16> CONF0_P<17> CONF0_P<18>
                           + CONF0_P<19> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4>
                           + CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8> CONF1_N<9> CONF1_N<10>
                           + CONF1_N<11> CONF1_N<12> CONF1_N<13> CONF1_N<14> CONF1_N<15> CONF1_N<16>
                           + CONF1_N<17> CONF1_N<18> CONF1_N<19> CONF1_P<0> CONF1_P<1> CONF1_P<2>
                           + CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8>
                           + CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12> CONF1_P<13> CONF1_P<14>
                           + CONF1_P<15> CONF1_P<16> CONF1_P<17> CONF1_P<18> CONF1_P<19> CONF_DEC<0>
                           + CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5> CONF_DEC<6>
                           + CONF_DEC<7> CONF_DEC<8> CONF_DEC<9> CONF_MAXCYCLES<0> CONF_MAXCYCLES<1>
                           + CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5>
                           + CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> CONF_WAITCYCLES<0>
                           + CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
                           + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                           + CONF_WAITCYCLES<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L FF<0>
                           + FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> FF<8> FF<9> RAND_OUT READY
                           + RST RST' VDD VSS
    Xi7 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_DEC<4> CONF_DEC<5> CONF_DEC<6>
        + CONF_DEC<7> CONF_DEC<8> CONF_DEC<9> FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> FF<8>
        + FF<9> RAND_OUT VDD VSS dec_10_conf_0
    Xi1 net35<0> net35<1> net35<2> net35<3> net35<4> BUF0_P<0> BUF0_P<1> BUF0_P<2> BUF0_P<3>
        + BUF0_P<4> net34<0> net34<1> net34<2> net34<3> net34<4> BUF1_P<0> BUF1_P<1> BUF1_P<2>
        + BUF1_P<3> BUF1_P<4> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_N<4> CONF0_N<5>
        + CONF0_N<6> CONF0_N<7> CONF0_N<8> CONF0_N<9> CONF0_N<10> CONF0_N<11> CONF0_N<12>
        + CONF0_N<13> CONF0_N<14> CONF0_N<15> CONF0_N<16> CONF0_N<17> CONF0_N<18> CONF0_N<19>
        + CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7>
        + CONF0_P<8> CONF0_P<9> CONF0_P<10> CONF0_P<11> CONF0_P<12> CONF0_P<13> CONF0_P<14>
        + CONF0_P<15> CONF0_P<16> CONF0_P<17> CONF0_P<18> CONF0_P<19> CONF1_N<0> CONF1_N<1>
        + CONF1_N<2> CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_N<8> CONF1_N<9>
        + CONF1_N<10> CONF1_N<11> CONF1_N<12> CONF1_N<13> CONF1_N<14> CONF1_N<15> CONF1_N<16>
        + CONF1_N<17> CONF1_N<18> CONF1_N<19> CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> CONF1_P<4>
        + CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF1_P<8> CONF1_P<9> CONF1_P<10> CONF1_P<11> CONF1_P<12>
        + CONF1_P<13> CONF1_P<14> CONF1_P<15> CONF1_P<16> CONF1_P<17> CONF1_P<18> CONF1_P<19>
        + EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> FF<8>
        + FF<9> RST RST' VDD VSS tdc_2e_4b_diff_np_4lin_buf
    Xi2 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
        + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7>
        + CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
        + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
        + FF<0> FF<1> FF<2> FF<3> FF<4> FF<5> FF<6> FF<7> FF<8> FF<9> BUF0_P<0> READY RST RST' VDD
        + VSS tdc_ready_6
.ENDS

.SUBCKT tdc_2e_1b_diff_np_4lin_buf BUF0_N<0> BUF0_N<1> BUF0_P<0> BUF0_P<1> BUF1_N<0> BUF1_N<1>
                                   + BUF1_P<0> BUF1_P<1> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
                                   + CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_P<0>
                                   + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5>
                                   + CONF0_P<6> CONF0_P<7> CONF1_N<0> CONF1_N<1> CONF1_N<2>
                                   + CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
                                   + CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> CONF1_P<4>
                                   + CONF1_P<5> CONF1_P<6> CONF1_P<7> EDGE0_N EDGE0_P EDGE1_N
                                   + EDGE1_P FF0<0> FF0<1> FF1<0> FF1<1> RST RST' VDD VSS
    Xi13 BUF0_N<1> BUF0_P<1> BUF1_N<1> BUF1_P<1> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7>
         + CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7>
         + CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> FF0<1> FF1<1> INT0_N<0> INT0_P<0> INT1_N<0>
         + INT1_P<0> NAND0<0> NAND0<1> NAND1<0> NAND1<1> INT0_N<1> INT0_P<1> INT1_N<1> INT1_P<1> RST
         + RST' VDD VSS tdc_2stage_diff_np_4lin_buf
    Xi12 BUF0_N<0> BUF0_P<0> BUF1_N<0> BUF1_P<0> CONF0_N<0> CONF0_N<1> CONF0_N<2> CONF0_N<3>
         + CONF0_P<0> CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3>
         + CONF1_P<0> CONF1_P<1> CONF1_P<2> CONF1_P<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P FF0<0> FF1<0>
         + INT1_N<1> INT1_P<1> INT0_N<1> INT0_P<1> NAND1<1> NAND0<0> NAND0<1> NAND1<0> INT0_N<0>
         + INT0_P<0> INT1_N<0> INT1_P<0> RST RST' VDD VSS tdc_2stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT dec_4_conf_0 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> FF_IN<0> FF_IN<1> FF_IN<2>
                     + FF_IN<3> RAND_OUT VDD VSS
    Xi27 CONF_DEC<3> FF_IN<3> FF_IN<2> STAGE<3> VDD VSS dec_stage
    Xi21 CONF_DEC<2> FF_IN<2> FF_IN<1> STAGE<2> VDD VSS dec_stage
    Xi19 CONF_DEC<1> FF_IN<1> FF_IN<0> STAGE<1> VDD VSS dec_stage
    Xi18 CONF_DEC<0> FF_IN<0> FF_IN<3> STAGE<0> VDD VSS dec_stage
    Xi26 net026 net023 RAND_OUT VDD VSS nor2
    Xi25 STAGE<2> STAGE<3> net023 VDD VSS nand2
    Xi24 STAGE<0> STAGE<1> net026 VDD VSS nand2
.ENDS

.SUBCKT ff_ready_2 FF0<0> FF0<1> FF1<0> FF1<1> FF_READY RST RST' VDD VSS
    Xi2 FF_NOR0 FF_NOR1 FF_NAND VDD VSS nand2
    Xi3 FF_NAND FF_READY net18 RST RST' VDD VSS dff_st_ar_dh
    Xi0 FF0<0> FF0<1> FF_NOR0 VDD VSS nor2
    Xi1 FF1<0> FF1<1> FF_NOR1 VDD VSS nor2
.ENDS

.SUBCKT tdc_ready_2 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
                    + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6>
                    + CONF_MAXCYCLES<7> CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2>
                    + CONF_WAITCYCLES<3> CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                    + CONF_WAITCYCLES<7> ENABLE_E2L FF0<0> FF0<1> FF1<0> FF1<1> INT READY RST RST'
                    + VDD VSS
    Xi20 CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4>
         + CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> INT net017 RST RST' VDD VSS
         + max_ready
    Xi32 ALARM<0> net19 net027 READY_I VDD VSS nand3
    Xi19 CLK CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
         + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
         + INT RST RST' VDD VSS WAIT_Ready wait_ready
    Xi28 WAIT_Ready net19 VDD VSS inv
    Xi27 FF_Ready ALARM<0> VDD VSS inv
    Xi30 READY_I READY Ready' RST RST' VDD VSS dff_st_ar_dh
    Xi33 net017 Ready' ALARM<1> net027 RST RST' VDD VSS dff_st_ar
    Xi18 FF0<0> FF0<1> FF1<0> FF1<1> FF_Ready RST RST' VDD VSS ff_ready_2
.ENDS

.SUBCKT tdc_1b_diff_branch ALARM<0> ALARM<1> BUF1_P<0> CLK CONF0_N<0> CONF0_N<1> CONF0_N<2>
                           + CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_P<0>
                           + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6>
                           + CONF0_P<7> CONF1_N<0> CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4>
                           + CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_P<0> CONF1_P<1> CONF1_P<2>
                           + CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> CONF_DEC<0>
                           + CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> CONF_MAXCYCLES<0> CONF_MAXCYCLES<1>
                           + CONF_MAXCYCLES<2> CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5>
                           + CONF_MAXCYCLES<6> CONF_MAXCYCLES<7> CONF_WAITCYCLES<0>
                           + CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
                           + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6>
                           + CONF_WAITCYCLES<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L FF<0>
                           + FF<1> FF<2> FF<3> RAND_OUT READY RST RST' VDD VSS
    Xi1 net31<0> net31<1> BUF0_P<0> BUF0_P<1> net30<0> net30<1> BUF1_P<0> BUF1_P<1> CONF0_N<0>
        + CONF0_N<1> CONF0_N<2> CONF0_N<3> CONF0_N<4> CONF0_N<5> CONF0_N<6> CONF0_N<7> CONF0_P<0>
        + CONF0_P<1> CONF0_P<2> CONF0_P<3> CONF0_P<4> CONF0_P<5> CONF0_P<6> CONF0_P<7> CONF1_N<0>
        + CONF1_N<1> CONF1_N<2> CONF1_N<3> CONF1_N<4> CONF1_N<5> CONF1_N<6> CONF1_N<7> CONF1_P<0>
        + CONF1_P<1> CONF1_P<2> CONF1_P<3> CONF1_P<4> CONF1_P<5> CONF1_P<6> CONF1_P<7> EDGE0_N
        + EDGE0_P EDGE1_N EDGE1_P FF<0> FF<1> FF<2> FF<3> RST RST' VDD VSS
        + tdc_2e_1b_diff_np_4lin_buf
    Xi7 CONF_DEC<0> CONF_DEC<1> CONF_DEC<2> CONF_DEC<3> FF<0> FF<1> FF<2> FF<3> RAND_OUT VDD VSS
        + dec_4_conf_0
    Xi2 ALARM<0> ALARM<1> CLK CONF_MAXCYCLES<0> CONF_MAXCYCLES<1> CONF_MAXCYCLES<2>
        + CONF_MAXCYCLES<3> CONF_MAXCYCLES<4> CONF_MAXCYCLES<5> CONF_MAXCYCLES<6> CONF_MAXCYCLES<7>
        + CONF_WAITCYCLES<0> CONF_WAITCYCLES<1> CONF_WAITCYCLES<2> CONF_WAITCYCLES<3>
        + CONF_WAITCYCLES<4> CONF_WAITCYCLES<5> CONF_WAITCYCLES<6> CONF_WAITCYCLES<7> ENABLE_E2L
        + FF<0> FF<1> FF<2> FF<3> BUF0_P<0> READY RST RST' VDD VSS tdc_ready_2
.ENDS

.SUBCKT trng_toplevel ALARM0<0> ALARM0<1> ALARM1<0> ALARM1<1> ALARM_DC CLK CONF_DEC0<0> CONF_DEC0<1>
                      + CONF_DEC0<2> CONF_DEC0<3> CONF_DEC0<4> CONF_DEC0<5> CONF_DEC0<6>
                      + CONF_DEC0<7> CONF_DEC0<8> CONF_DEC0<9> CONF_DEC1<0> CONF_DEC1<1>
                      + CONF_DEC1<2> CONF_DEC1<3> CONF_DEC1<4> CONF_DEC1<5> CONF_DEC1<6>
                      + CONF_DEC1<7> CONF_DEC1<8> CONF_DEC1<9> CONF_SELDC<0> CONF_SELDC<1>
                      + CONF_SELTDC<0> CONF_SELTDC<1> CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
                      + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7>
                      + CONF_TDC00N<8> CONF_TDC00N<9> CONF_TDC00N<10> CONF_TDC00N<11>
                      + CONF_TDC00N<12> CONF_TDC00N<13> CONF_TDC00N<14> CONF_TDC00N<15>
                      + CONF_TDC00N<16> CONF_TDC00N<17> CONF_TDC00N<18> CONF_TDC00N<19>
                      + CONF_TDC00P<0> CONF_TDC00P<1> CONF_TDC00P<2> CONF_TDC00P<3> CONF_TDC00P<4>
                      + CONF_TDC00P<5> CONF_TDC00P<6> CONF_TDC00P<7> CONF_TDC00P<8> CONF_TDC00P<9>
                      + CONF_TDC00P<10> CONF_TDC00P<11> CONF_TDC00P<12> CONF_TDC00P<13>
                      + CONF_TDC00P<14> CONF_TDC00P<15> CONF_TDC00P<16> CONF_TDC00P<17>
                      + CONF_TDC00P<18> CONF_TDC00P<19> CONF_TDC01N<0> CONF_TDC01N<1> CONF_TDC01N<2>
                      + CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5> CONF_TDC01N<6> CONF_TDC01N<7>
                      + CONF_TDC01N<8> CONF_TDC01N<9> CONF_TDC01N<10> CONF_TDC01N<11>
                      + CONF_TDC01N<12> CONF_TDC01N<13> CONF_TDC01N<14> CONF_TDC01N<15>
                      + CONF_TDC01N<16> CONF_TDC01N<17> CONF_TDC01N<18> CONF_TDC01N<19>
                      + CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2> CONF_TDC01P<3> CONF_TDC01P<4>
                      + CONF_TDC01P<5> CONF_TDC01P<6> CONF_TDC01P<7> CONF_TDC01P<8> CONF_TDC01P<9>
                      + CONF_TDC01P<10> CONF_TDC01P<11> CONF_TDC01P<12> CONF_TDC01P<13>
                      + CONF_TDC01P<14> CONF_TDC01P<15> CONF_TDC01P<16> CONF_TDC01P<17>
                      + CONF_TDC01P<18> CONF_TDC01P<19> CONF_TDC4B CONF_TDC10N<0> CONF_TDC10N<1>
                      + CONF_TDC10N<2> CONF_TDC10N<3> CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6>
                      + CONF_TDC10N<7> CONF_TDC10N<8> CONF_TDC10N<9> CONF_TDC10N<10> CONF_TDC10N<11>
                      + CONF_TDC10N<12> CONF_TDC10N<13> CONF_TDC10N<14> CONF_TDC10N<15>
                      + CONF_TDC10N<16> CONF_TDC10N<17> CONF_TDC10N<18> CONF_TDC10N<19>
                      + CONF_TDC10P<0> CONF_TDC10P<1> CONF_TDC10P<2> CONF_TDC10P<3> CONF_TDC10P<4>
                      + CONF_TDC10P<5> CONF_TDC10P<6> CONF_TDC10P<7> CONF_TDC10P<8> CONF_TDC10P<9>
                      + CONF_TDC10P<10> CONF_TDC10P<11> CONF_TDC10P<12> CONF_TDC10P<13>
                      + CONF_TDC10P<14> CONF_TDC10P<15> CONF_TDC10P<16> CONF_TDC10P<17>
                      + CONF_TDC10P<18> CONF_TDC10P<19> CONF_TDC11N<0> CONF_TDC11N<1> CONF_TDC11N<2>
                      + CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5> CONF_TDC11N<6> CONF_TDC11N<7>
                      + CONF_TDC11N<8> CONF_TDC11N<9> CONF_TDC11N<10> CONF_TDC11N<11>
                      + CONF_TDC11N<12> CONF_TDC11N<13> CONF_TDC11N<14> CONF_TDC11N<15>
                      + CONF_TDC11N<16> CONF_TDC11N<17> CONF_TDC11N<18> CONF_TDC11N<19>
                      + CONF_TDC11P<0> CONF_TDC11P<1> CONF_TDC11P<2> CONF_TDC11P<3> CONF_TDC11P<4>
                      + CONF_TDC11P<5> CONF_TDC11P<6> CONF_TDC11P<7> CONF_TDC11P<8> CONF_TDC11P<9>
                      + CONF_TDC11P<10> CONF_TDC11P<11> CONF_TDC11P<12> CONF_TDC11P<13>
                      + CONF_TDC11P<14> CONF_TDC11P<15> CONF_TDC11P<16> CONF_TDC11P<17>
                      + CONF_TDC11P<18> CONF_TDC11P<19> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2>
                      + CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
                      + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3>
                      + CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> DCEDGE0<1>
                      + DCEDGE0<2> DCEDGE0<3> DCEDGE1<1> DCEDGE1<2> DCEDGE1<3> DCEDGE2<1> DCEDGE2<2>
                      + DCEDGE2<3> ENABLE_E2L ENABLE_MERO FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF0<5>
                      + FF0<6> FF0<7> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF1<5> FF1<6> FF1<7> INT0
                      + INT1 MERO_INT<0> MERO_INT<1> MERO_INT<2> RAND_OUT0 RAND_OUT1 READY0 READY1
                      + RST RST' SEL_DCEDGE<0> SEL_DCEDGE<1> TDC0_FF4<0> TDC0_FF5<0> TDC0_FF5<3>
                      + TDC0_FF6<0> TDC0_FF6<1> TDC0_FF6<3> TDC0_FF7<0> TDC0_FF7<1> TDC0_FF7<3>
                      + TDC1_FF4<0> TDC1_FF5<0> TDC1_FF5<3> TDC1_FF6<0> TDC1_FF6<1> TDC1_FF6<3>
                      + TDC1_FF7<0> TDC1_FF7<1> TDC1_FF7<3> VDD_CORE VDD_DC VDD_TDC VSS
    Xi81 TDC03_FF<0> TDC03_FF<1> TDC03_FF<2> TDC03_FF<3> TDC03_FF<4> TDC03_FF<5> TDC03_FF<6>
         + TDC03_FF<7> TDC03_FF<8> TDC03_FF<9> TDC13_FF<0> TDC13_FF<1> TDC13_FF<2> TDC13_FF<3>
         + TDC13_FF<4> TDC13_FF<5> TDC13_FF<6> TDC13_FF<7> TDC13_FF<8> TDC13_FF<9> TDC0_FF0<3>
         + TDC0_FF1<3> TDC0_FF2<3> TDC0_FF3<3> TDC0_FF4<3> TDC1_FF0<3> TDC1_FF1<3> TDC1_FF2<3>
         + TDC1_FF3<3> TDC1_FF4<3> CONF_TDC4B VDD_CORE VSS mux2_10x
    Xi77 TDC1_ALARM0<1> TDC1_ALARM1<1> TDC1_INT<1> CLK CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2>
         + CONF_TDC10N<3> CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10N<8>
         + CONF_TDC10N<9> CONF_TDC10N<10> CONF_TDC10N<11> CONF_TDC10P<0> CONF_TDC10P<1>
         + CONF_TDC10P<2> CONF_TDC10P<3> CONF_TDC10P<4> CONF_TDC10P<5> CONF_TDC10P<6> CONF_TDC10P<7>
         + CONF_TDC10P<8> CONF_TDC10P<9> CONF_TDC10P<10> CONF_TDC10P<11> CONF_TDC11N<0>
         + CONF_TDC11N<1> CONF_TDC11N<2> CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5> CONF_TDC11N<6>
         + CONF_TDC11N<7> CONF_TDC11N<8> CONF_TDC11N<9> CONF_TDC11N<10> CONF_TDC11N<11>
         + CONF_TDC11P<0> CONF_TDC11P<1> CONF_TDC11P<2> CONF_TDC11P<3> CONF_TDC11P<4> CONF_TDC11P<5>
         + CONF_TDC11P<6> CONF_TDC11P<7> CONF_TDC11P<8> CONF_TDC11P<9> CONF_TDC11P<10>
         + CONF_TDC11P<11> CONF_DEC1<0> CONF_DEC1<1> CONF_DEC1<2> CONF_DEC1<3> CONF_DEC1<4>
         + CONF_DEC1<5> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4>
         + CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7> CONF_TDCWAIT<0> CONF_TDCWAIT<1>
         + CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6>
         + CONF_TDCWAIT<7> EDGE1_N EDGE1_P EDGE2_N EDGE2_P ENABLE_E2L TDC1_FF0<1> TDC1_FF1<1>
         + TDC1_FF2<1> TDC1_FF3<1> TDC1_FF4<1> TDC1_FF5<1> TDC1_RANDOUT<1> TDC1_READY<1> RST RST'
         + VDD_TDC_INT1<1> VSS tdc_2b_diff_branch
    Xi73 TDC0_ALARM0<1> TDC0_ALARM1<1> TDC0_INT<1> CLK CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
         + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7> CONF_TDC00N<8>
         + CONF_TDC00N<9> CONF_TDC00N<10> CONF_TDC00N<11> CONF_TDC00P<0> CONF_TDC00P<1>
         + CONF_TDC00P<2> CONF_TDC00P<3> CONF_TDC00P<4> CONF_TDC00P<5> CONF_TDC00P<6> CONF_TDC00P<7>
         + CONF_TDC00P<8> CONF_TDC00P<9> CONF_TDC00P<10> CONF_TDC00P<11> CONF_TDC01N<0>
         + CONF_TDC01N<1> CONF_TDC01N<2> CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5> CONF_TDC01N<6>
         + CONF_TDC01N<7> CONF_TDC01N<8> CONF_TDC01N<9> CONF_TDC01N<10> CONF_TDC01N<11>
         + CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2> CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5>
         + CONF_TDC01P<6> CONF_TDC01P<7> CONF_TDC01P<8> CONF_TDC01P<9> CONF_TDC01P<10>
         + CONF_TDC01P<11> CONF_DEC0<0> CONF_DEC0<1> CONF_DEC0<2> CONF_DEC0<3> CONF_DEC0<4>
         + CONF_DEC0<5> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4>
         + CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7> CONF_TDCWAIT<0> CONF_TDCWAIT<1>
         + CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6>
         + CONF_TDCWAIT<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L TDC0_FF0<1> TDC0_FF1<1>
         + TDC0_FF2<1> TDC0_FF3<1> TDC0_FF4<1> TDC0_FF5<1> TDC0_RANDOUT<1> TDC0_READY<1> RST RST'
         + VDD_TDC_INT0<1> VSS tdc_2b_diff_branch
    Xi78 TDC1_ALARM0<2> TDC1_ALARM1<2> TDC1_INT<2> CLK CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2>
         + CONF_TDC10N<3> CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10N<8>
         + CONF_TDC10N<9> CONF_TDC10N<10> CONF_TDC10N<11> CONF_TDC10N<12> CONF_TDC10N<13>
         + CONF_TDC10N<14> CONF_TDC10N<15> CONF_TDC10P<0> CONF_TDC10P<1> CONF_TDC10P<2>
         + CONF_TDC10P<3> CONF_TDC10P<4> CONF_TDC10P<5> CONF_TDC10P<6> CONF_TDC10P<7> CONF_TDC10P<8>
         + CONF_TDC10P<9> CONF_TDC10P<10> CONF_TDC10P<11> CONF_TDC10P<12> CONF_TDC10P<13>
         + CONF_TDC10P<14> CONF_TDC10P<15> CONF_TDC11N<0> CONF_TDC11N<1> CONF_TDC11N<2>
         + CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5> CONF_TDC11N<6> CONF_TDC11N<7> CONF_TDC11N<8>
         + CONF_TDC11N<9> CONF_TDC11N<10> CONF_TDC11N<11> CONF_TDC11N<12> CONF_TDC11N<13>
         + CONF_TDC11N<14> CONF_TDC11N<15> CONF_TDC11P<0> CONF_TDC11P<1> CONF_TDC11P<2>
         + CONF_TDC11P<3> CONF_TDC11P<4> CONF_TDC11P<5> CONF_TDC11P<6> CONF_TDC11P<7> CONF_TDC11P<8>
         + CONF_TDC11P<9> CONF_TDC11P<10> CONF_TDC11P<11> CONF_TDC11P<12> CONF_TDC11P<13>
         + CONF_TDC11P<14> CONF_TDC11P<15> CONF_DEC1<0> CONF_DEC1<1> CONF_DEC1<2> CONF_DEC1<3>
         + CONF_DEC1<4> CONF_DEC1<5> CONF_DEC1<6> CONF_DEC1<7> CONF_TDCMAX<0> CONF_TDCMAX<1>
         + CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
         + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4>
         + CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> EDGE1_N EDGE1_P EDGE2_N EDGE2_P
         + ENABLE_E2L TDC1_FF0<2> TDC1_FF1<2> TDC1_FF2<2> TDC1_FF3<2> TDC1_FF4<2> TDC1_FF5<2>
         + TDC1_FF6<2> TDC1_FF7<2> TDC1_RANDOUT<2> TDC1_READY<2> RST RST' VDD_TDC_INT1<2> VSS
         + tdc_3b_diff_branch
    Xi74 TDC0_ALARM0<2> TDC0_ALARM1<2> TDC0_INT<2> CLK CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
         + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7> CONF_TDC00N<8>
         + CONF_TDC00N<9> CONF_TDC00N<10> CONF_TDC00N<11> CONF_TDC00N<12> CONF_TDC00N<13>
         + CONF_TDC00N<14> CONF_TDC00N<15> CONF_TDC00P<0> CONF_TDC00P<1> CONF_TDC00P<2>
         + CONF_TDC00P<3> CONF_TDC00P<4> CONF_TDC00P<5> CONF_TDC00P<6> CONF_TDC00P<7> CONF_TDC00P<8>
         + CONF_TDC00P<9> CONF_TDC00P<10> CONF_TDC00P<11> CONF_TDC00P<12> CONF_TDC00P<13>
         + CONF_TDC00P<14> CONF_TDC00P<15> CONF_TDC01N<0> CONF_TDC01N<1> CONF_TDC01N<2>
         + CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5> CONF_TDC01N<6> CONF_TDC01N<7> CONF_TDC01N<8>
         + CONF_TDC01N<9> CONF_TDC01N<10> CONF_TDC01N<11> CONF_TDC01N<12> CONF_TDC01N<13>
         + CONF_TDC01N<14> CONF_TDC01N<15> CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2>
         + CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5> CONF_TDC01P<6> CONF_TDC01P<7> CONF_TDC01P<8>
         + CONF_TDC01P<9> CONF_TDC01P<10> CONF_TDC01P<11> CONF_TDC01P<12> CONF_TDC01P<13>
         + CONF_TDC01P<14> CONF_TDC01P<15> CONF_DEC0<0> CONF_DEC0<1> CONF_DEC0<2> CONF_DEC0<3>
         + CONF_DEC0<4> CONF_DEC0<5> CONF_DEC0<6> CONF_DEC0<7> CONF_TDCMAX<0> CONF_TDCMAX<1>
         + CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
         + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4>
         + CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P
         + ENABLE_E2L TDC0_FF0<2> TDC0_FF1<2> TDC0_FF2<2> TDC0_FF3<2> TDC0_FF4<2> TDC0_FF5<2>
         + TDC0_FF6<2> TDC0_FF7<2> TDC0_RANDOUT<2> TDC0_READY<2> RST RST' VDD_TDC_INT0<2> VSS
         + tdc_3b_diff_branch
    Xi80 ALARM_DC CONF_SELDC<0> CONF_SELDC<1> DCEDGE0<1> DCEDGE0<2> DCEDGE0<3> DCEDGE1<1> DCEDGE1<2>
         + DCEDGE1<3> DCEDGE2<1> DCEDGE2<2> DCEDGE2<3> EDGE0_N EDGE0_P EDGE1_N EDGE1_P EDGE2_N
         + EDGE2_P ENABLE_E2L ENABLE_MERO MERO_INT<0> MERO_INT<1> MERO_INT<2> RST RST' SEL_DCEDGE<0>
         + SEL_DCEDGE<1> VDD_CORE VDD_DC VSS dc_collection
    Xi56 TDC1_FF7<0> TDC1_FF7<1> TDC1_FF7<2> TDC1_FF7<3> FF1<7> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi55 TDC1_FF6<0> TDC1_FF6<1> TDC1_FF6<2> TDC1_FF6<3> FF1<6> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi54 TDC1_FF5<0> TDC1_FF5<1> TDC1_FF5<2> TDC1_FF5<3> FF1<5> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi53 TDC1_FF4<0> TDC1_FF4<1> TDC1_FF4<2> TDC1_FF4<3> FF1<4> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi52 TDC1_FF3<0> TDC1_FF3<1> TDC1_FF3<2> TDC1_FF3<3> FF1<3> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi51 TDC1_FF2<0> TDC1_FF2<1> TDC1_FF2<2> TDC1_FF2<3> FF1<2> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi50 TDC1_FF1<0> TDC1_FF1<1> TDC1_FF1<2> TDC1_FF1<3> FF1<1> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi49 TDC0_FF7<0> TDC0_FF7<1> TDC0_FF7<2> TDC0_FF7<3> FF0<7> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi48 TDC0_FF6<0> TDC0_FF6<1> TDC0_FF6<2> TDC0_FF6<3> FF0<6> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi47 TDC0_FF5<0> TDC0_FF5<1> TDC0_FF5<2> TDC0_FF5<3> FF0<5> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi46 TDC0_FF4<0> TDC0_FF4<1> TDC0_FF4<2> TDC0_FF4<3> FF0<4> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi45 TDC0_FF3<0> TDC0_FF3<1> TDC0_FF3<2> TDC0_FF3<3> FF0<3> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi44 TDC0_FF2<0> TDC0_FF2<1> TDC0_FF2<2> TDC0_FF2<3> FF0<2> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi43 TDC0_FF1<0> TDC0_FF1<1> TDC0_FF1<2> TDC0_FF1<3> FF0<1> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi42 TDC1_RANDOUT<0> TDC1_RANDOUT<1> TDC1_RANDOUT<2> TDC1_RANDOUT<3> RAND_OUT1 CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi41 TDC1_FF0<0> TDC1_FF0<1> TDC1_FF0<2> TDC1_FF0<3> FF1<0> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi40 TDC1_ALARM1<0> TDC1_ALARM1<1> TDC1_ALARM1<2> TDC1_ALARM1<3> ALARM1<1> CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi39 TDC1_ALARM0<0> TDC1_ALARM0<1> TDC1_ALARM0<2> TDC1_ALARM0<3> ALARM1<0> CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi38 TDC1_INT<0> TDC1_INT<1> TDC1_INT<2> TDC1_INT<3> INT1 CONF_SELTDC<0> CONF_SELTDC<1> VDD_CORE
         + VSS mux4
    Xi37 TDC1_READY<0> TDC1_READY<1> TDC1_READY<2> TDC1_READY<3> READY1 CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi36 TDC0_FF0<0> TDC0_FF0<1> TDC0_FF0<2> TDC0_FF0<3> FF0<0> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS mux4
    Xi35 TDC0_ALARM1<0> TDC0_ALARM1<1> TDC0_ALARM1<2> TDC0_ALARM1<3> ALARM0<1> CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi34 TDC0_ALARM0<0> TDC0_ALARM0<1> TDC0_ALARM0<2> TDC0_ALARM0<3> ALARM0<0> CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi33 TDC0_INT<0> TDC0_INT<1> TDC0_INT<2> TDC0_INT<3> INT0 CONF_SELTDC<0> CONF_SELTDC<1> VDD_CORE
         + VSS mux4
    Xi32 TDC0_READY<0> TDC0_READY<1> TDC0_READY<2> TDC0_READY<3> READY0 CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi31 TDC0_RANDOUT<0> TDC0_RANDOUT<1> TDC0_RANDOUT<2> TDC0_RANDOUT<3> RAND_OUT0 CONF_SELTDC<0>
         + CONF_SELTDC<1> VDD_CORE VSS mux4
    Xi69 SELTDC_DEC<3> VDD_TDC VDD_TDC_INT1<3> VSS vdd_gate_1ma
    Xi68 SELTDC_DEC<3> VDD_TDC VDD_TDC_INT0<3> VSS vdd_gate_1ma
    Xi67 SELTDC_DEC<2> VDD_TDC VDD_TDC_INT0<2> VSS vdd_gate_1ma
    Xi66 SELTDC_DEC<2> VDD_TDC VDD_TDC_INT1<2> VSS vdd_gate_1ma
    Xi63 SELTDC_DEC<1> VDD_TDC VDD_TDC_INT0<1> VSS vdd_gate_1ma
    Xi62 SELTDC_DEC<1> VDD_TDC VDD_TDC_INT1<1> VSS vdd_gate_1ma
    Xi58 SELTDC_DEC<0> VDD_TDC VDD_TDC_INT1<0> VSS vdd_gate_1ma
    Xi57 SELTDC_DEC<0> VDD_TDC VDD_TDC_INT0<0> VSS vdd_gate_1ma
    Xi59 SELTDC_DEC<0> SELTDC_DEC<1> SELTDC_DEC<2> SELTDC_DEC<3> CONF_SELTDC<0> CONF_SELTDC<1>
         + VDD_CORE VSS dec4_inverted
    Xi75 TDC0_ALARM0<3> TDC0_ALARM1<3> TDC0_INT<3> CLK CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
         + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7> CONF_TDC00N<8>
         + CONF_TDC00N<9> CONF_TDC00N<10> CONF_TDC00N<11> CONF_TDC00N<12> CONF_TDC00N<13>
         + CONF_TDC00N<14> CONF_TDC00N<15> CONF_TDC00N<16> CONF_TDC00N<17> CONF_TDC00N<18>
         + CONF_TDC00N<19> CONF_TDC00P<0> CONF_TDC00P<1> CONF_TDC00P<2> CONF_TDC00P<3>
         + CONF_TDC00P<4> CONF_TDC00P<5> CONF_TDC00P<6> CONF_TDC00P<7> CONF_TDC00P<8> CONF_TDC00P<9>
         + CONF_TDC00P<10> CONF_TDC00P<11> CONF_TDC00P<12> CONF_TDC00P<13> CONF_TDC00P<14>
         + CONF_TDC00P<15> CONF_TDC00P<16> CONF_TDC00P<17> CONF_TDC00P<18> CONF_TDC00P<19>
         + CONF_TDC01N<0> CONF_TDC01N<1> CONF_TDC01N<2> CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5>
         + CONF_TDC01N<6> CONF_TDC01N<7> CONF_TDC01N<8> CONF_TDC01N<9> CONF_TDC01N<10>
         + CONF_TDC01N<11> CONF_TDC01N<12> CONF_TDC01N<13> CONF_TDC01N<14> CONF_TDC01N<15>
         + CONF_TDC01N<16> CONF_TDC01N<17> CONF_TDC01N<18> CONF_TDC01N<19> CONF_TDC01P<0>
         + CONF_TDC01P<1> CONF_TDC01P<2> CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5> CONF_TDC01P<6>
         + CONF_TDC01P<7> CONF_TDC01P<8> CONF_TDC01P<9> CONF_TDC01P<10> CONF_TDC01P<11>
         + CONF_TDC01P<12> CONF_TDC01P<13> CONF_TDC01P<14> CONF_TDC01P<15> CONF_TDC01P<16>
         + CONF_TDC01P<17> CONF_TDC01P<18> CONF_TDC01P<19> CONF_DEC0<0> CONF_DEC0<1> CONF_DEC0<2>
         + CONF_DEC0<3> CONF_DEC0<4> CONF_DEC0<5> CONF_DEC0<6> CONF_DEC0<7> CONF_DEC0<8>
         + CONF_DEC0<9> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4>
         + CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7> CONF_TDCWAIT<0> CONF_TDCWAIT<1>
         + CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6>
         + CONF_TDCWAIT<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P ENABLE_E2L TDC03_FF<0> TDC03_FF<1>
         + TDC03_FF<2> TDC03_FF<3> TDC03_FF<4> TDC03_FF<5> TDC03_FF<6> TDC03_FF<7> TDC03_FF<8>
         + TDC03_FF<9> TDC0_RANDOUT<3> TDC0_READY<3> RST RST' VDD_TDC_INT0<3> VSS tdc_4b_diff_branch
    Xi79 TDC1_ALARM0<3> TDC1_ALARM1<3> TDC1_INT<3> CLK CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2>
         + CONF_TDC10N<3> CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10N<8>
         + CONF_TDC10N<9> CONF_TDC10N<10> CONF_TDC10N<11> CONF_TDC10N<12> CONF_TDC10N<13>
         + CONF_TDC10N<14> CONF_TDC10N<15> CONF_TDC10N<16> CONF_TDC10N<17> CONF_TDC10N<18>
         + CONF_TDC10N<19> CONF_TDC10P<0> CONF_TDC10P<1> CONF_TDC10P<2> CONF_TDC10P<3>
         + CONF_TDC10P<4> CONF_TDC10P<5> CONF_TDC10P<6> CONF_TDC10P<7> CONF_TDC10P<8> CONF_TDC10P<9>
         + CONF_TDC10P<10> CONF_TDC10P<11> CONF_TDC10P<12> CONF_TDC10P<13> CONF_TDC10P<14>
         + CONF_TDC10P<15> CONF_TDC10P<16> CONF_TDC10P<17> CONF_TDC10P<18> CONF_TDC10P<19>
         + CONF_TDC11N<0> CONF_TDC11N<1> CONF_TDC11N<2> CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5>
         + CONF_TDC11N<6> CONF_TDC11N<7> CONF_TDC11N<8> CONF_TDC11N<9> CONF_TDC11N<10>
         + CONF_TDC11N<11> CONF_TDC11N<12> CONF_TDC11N<13> CONF_TDC11N<14> CONF_TDC11N<15>
         + CONF_TDC11N<16> CONF_TDC11N<17> CONF_TDC11N<18> CONF_TDC11N<19> CONF_TDC11P<0>
         + CONF_TDC11P<1> CONF_TDC11P<2> CONF_TDC11P<3> CONF_TDC11P<4> CONF_TDC11P<5> CONF_TDC11P<6>
         + CONF_TDC11P<7> CONF_TDC11P<8> CONF_TDC11P<9> CONF_TDC11P<10> CONF_TDC11P<11>
         + CONF_TDC11P<12> CONF_TDC11P<13> CONF_TDC11P<14> CONF_TDC11P<15> CONF_TDC11P<16>
         + CONF_TDC11P<17> CONF_TDC11P<18> CONF_TDC11P<19> CONF_DEC1<0> CONF_DEC1<1> CONF_DEC1<2>
         + CONF_DEC1<3> CONF_DEC1<4> CONF_DEC1<5> CONF_DEC1<6> CONF_DEC1<7> CONF_DEC1<8>
         + CONF_DEC1<9> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2> CONF_TDCMAX<3> CONF_TDCMAX<4>
         + CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7> CONF_TDCWAIT<0> CONF_TDCWAIT<1>
         + CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6>
         + CONF_TDCWAIT<7> EDGE1_N EDGE1_P EDGE2_N EDGE2_P ENABLE_E2L TDC13_FF<0> TDC13_FF<1>
         + TDC13_FF<2> TDC13_FF<3> TDC13_FF<4> TDC13_FF<5> TDC13_FF<6> TDC13_FF<7> TDC13_FF<8>
         + TDC13_FF<9> TDC1_RANDOUT<3> TDC1_READY<3> RST RST' VDD_TDC_INT1<3> VSS tdc_4b_diff_branch
    Xi72 TDC0_ALARM0<0> TDC0_ALARM1<0> TDC0_INT<0> CLK CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
         + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7> CONF_TDC00P<0>
         + CONF_TDC00P<1> CONF_TDC00P<2> CONF_TDC00P<3> CONF_TDC00P<4> CONF_TDC00P<5> CONF_TDC00P<6>
         + CONF_TDC00P<7> CONF_TDC01N<0> CONF_TDC01N<1> CONF_TDC01N<2> CONF_TDC01N<3> CONF_TDC01N<4>
         + CONF_TDC01N<5> CONF_TDC01N<6> CONF_TDC01N<7> CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2>
         + CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5> CONF_TDC01P<6> CONF_TDC01P<7> CONF_DEC0<0>
         + CONF_DEC0<1> CONF_DEC0<2> CONF_DEC0<3> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2>
         + CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
         + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4>
         + CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> EDGE0_N EDGE0_P EDGE1_N EDGE1_P
         + ENABLE_E2L TDC0_FF0<0> TDC0_FF1<0> TDC0_FF2<0> TDC0_FF3<0> TDC0_RANDOUT<0> TDC0_READY<0>
         + RST RST' VDD_TDC_INT0<0> VSS tdc_1b_diff_branch
    Xi76 TDC1_ALARM0<0> TDC1_ALARM1<0> TDC1_INT<0> CLK CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2>
         + CONF_TDC10N<3> CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10P<0>
         + CONF_TDC10P<1> CONF_TDC10P<2> CONF_TDC10P<3> CONF_TDC10P<4> CONF_TDC10P<5> CONF_TDC10P<6>
         + CONF_TDC10P<7> CONF_TDC11N<0> CONF_TDC11N<1> CONF_TDC11N<2> CONF_TDC11N<3> CONF_TDC11N<4>
         + CONF_TDC11N<5> CONF_TDC11N<6> CONF_TDC11N<7> CONF_TDC11P<0> CONF_TDC11P<1> CONF_TDC11P<2>
         + CONF_TDC11P<3> CONF_TDC11P<4> CONF_TDC11P<5> CONF_TDC11P<6> CONF_TDC11P<7> CONF_DEC1<0>
         + CONF_DEC1<1> CONF_DEC1<2> CONF_DEC1<3> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2>
         + CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
         + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4>
         + CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> EDGE1_N EDGE1_P EDGE2_N EDGE2_P
         + ENABLE_E2L TDC1_FF0<0> TDC1_FF1<0> TDC1_FF2<0> TDC1_FF3<0> TDC1_RANDOUT<0> TDC1_READY<0>
         + RST RST' VDD_TDC_INT1<0> VSS tdc_1b_diff_branch
.ENDS

.SUBCKT conf_control CAL_EN CAL_RO_EN CLK CTRL_RST DATA_READY RST RST' SER_READY STATE<0> STATE<1>
                     + STATE<2> STA_READY TDC_READY VDD VSS
    Xi2 CLK NEXTSTATE<2> STATE<2> STATE'<2> RST RST' VDD VSS dff_st_ar
    Xi1 CLK NEXTSTATE<1> STATE<1> STATE'<1> RST RST' VDD VSS dff_st_ar
    Xi0 CLK NEXTSTATE<0> STATE<0> STATE'<0> RST RST' VDD VSS dff_st_ar
    Xi14 STATE0_INT<0> STATE0_INT<1> STATE0_INT<2> STATE0_INT<3> NEXTSTATE<0> VDD VSS nand4
    Xi30 STATE'<0> STATE<1> STATE<2> net037 VDD VSS nand3
    Xi28 STATE<0> STATE'<1> STATE<2> net038 VDD VSS nand3
    Xi42 STATE'<0> STATE<1> STATE<2> STATE2_INT<2> VDD VSS nand3
    Xi23 STATE'<0> STATE<1> STA_READY STATE2_INT<1> VDD VSS nand3
    Xi43 STATE2_INT<0> STATE2_INT<1> STATE2_INT<2> NEXTSTATE<2> VDD VSS nand3
    Xi11 STATE<0> STATE<2> SER_READY' STATE0_INT<1> VDD VSS nand3
    Xi12 STATE<0> STATE<1> STATE<2> STATE0_INT<2> VDD VSS nand3
    Xi38 STATE<1> STATE<2> TDC_READY STATE0_INT<3> VDD VSS nand3
    Xi33 net044 CAL_RO_EN_I VDD VSS inv
    Xi31 net037 CAL_EN_I VDD VSS inv
    Xi29 net038 DATA_READY_I VDD VSS inv
    Xi45 SER_READY SER_READY' VDD VSS inv
    Xi32 STATE'<0> STATE<1> net044 VDD VSS nand2
    Xi34 CTRL_RST_INT<0> CTRL_RST_INT<1> CTRL_RST VDD VSS nand2
    Xi36 STATE'<1> STATE'<2> CTRL_RST_INT<0> VDD VSS nand2
    Xi22 STATE<0> STATE<2> STATE2_INT<0> VDD VSS nand2
    Xi41 STATE1_INT<0> STATE1_INT<1> NEXTSTATE<1> VDD VSS nand2
    Xi40 STATE<0> STATE'<2> STATE1_INT<1> VDD VSS nand2
    Xi39 STATE'<0> STATE<1> STATE1_INT<0> VDD VSS nand2
    Xi10 STATE'<1> STATE'<2> STATE0_INT<0> VDD VSS nand2
    Xi44 STATE<0> STATE'<2> CTRL_RST_INT<1> VDD VSS nand2
    Xi48 DATA_READY_I DATA_READY VDD VSS buffer
    Xi49 CAL_EN_I CAL_EN VDD VSS buffer
    Xi46 CAL_RO_EN_I CAL_RO_EN VDD VSS buffer
.ENDS

.SUBCKT asynccounter_16 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                        + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> Q' RST RST' VDD VSS
    Xi1 net12 OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> Q' RST RST' VDD VSS
        + asynccounter_8
    Xi0 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> net12 RST RST' VDD VSS
        + asynccounter_8
.ENDS

.SUBCKT inv_conf CONF'<0> CONF'<1> CONF'<2> CONF'<3> CONF<0> CONF<1> CONF<2> CONF<3> IN OUT VDD VSS
    Mm16 OUT IN VDD VDD p_mos l=60n w=120.0n m=1
    Mm7 OUT IN net16 VDD p_mos l=60n w=120.0n m=1
    Mm6 OUT IN net17 VDD p_mos l=60n w=120.0n m=1
    Mm5 OUT IN net18 VDD p_mos l=60n w=120.0n m=1
    Mm4 OUT IN net19 VDD p_mos l=60n w=120.0n m=1
    Mm3 net16 CONF'<3> VDD VDD p_mos l=60n w=120.0n m=1
    Mm2 net17 CONF'<2> VDD VDD p_mos l=60n w=120.0n m=1
    Mm1 net18 CONF'<1> VDD VDD p_mos l=60n w=120.0n m=1
    Mm0 net19 CONF'<0> VDD VDD p_mos l=60n w=120.0n m=1
    Mm17 OUT IN VSS VSS n_mos l=60n w=120.0n m=1
    Mm15 net20 CONF<3> VSS VSS n_mos l=60n w=120.0n m=1
    Mm14 OUT IN net20 VSS n_mos l=60n w=120.0n m=1
    Mm13 net21 CONF<2> VSS VSS n_mos l=60n w=120.0n m=1
    Mm12 OUT IN net21 VSS n_mos l=60n w=120.0n m=1
    Mm11 net22 CONF<1> VSS VSS n_mos l=60n w=120.0n m=1
    Mm10 OUT IN net22 VSS n_mos l=60n w=120.0n m=1
    Mm9 net23 CONF<0> VSS VSS n_mos l=60n w=120.0n m=1
    Mm8 OUT IN net23 VSS n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT ro_2i CONF'<0> CONF'<1> CONF'<2> CONF'<3> CONF'<4> CONF'<5> CONF'<6> CONF'<7> CONF<0>
              + CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> ENABLE OUT VDD VSS
    Xi1 CONF'<4> CONF'<5> CONF'<6> CONF'<7> CONF<4> CONF<5> CONF<6> CONF<7> INT OUT VDD VSS inv_conf
    Xi0 CONF'<0> CONF'<1> CONF'<2> CONF'<3> CONF<0> CONF<1> CONF<2> CONF<3> NAND_OUT INT VDD VSS
        + inv_conf
    Xi2 OUT ENABLE NAND_OUT VDD VSS nand2
.ENDS

.SUBCKT freqscaler3 CLK OUT<0> OUT<1> OUT<2> RST RST' VDD VSS
    Xi2 INT<1> OUT<2> net16 RST RST' VDD VSS tff_st_ar
    Xi1 INT<0> OUT<1> INT<1> RST RST' VDD VSS tff_st_ar
    Xi0 CLK OUT<0> INT<0> RST RST' VDD VSS tff_st_ar
.ENDS

.SUBCKT inv_sd IN OUT VDD VSS
    Mm0 OUT IN VSS VSS n_mos l=60n w=480.0n m=1
    Mm1 OUT IN VDD VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT inv_bank_8 IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> OUT<0> OUT<1> OUT<2> OUT<3>
                   + OUT<4> OUT<5> OUT<6> OUT<7> VDD VSS
    Xi7 IN<7> OUT<7> VDD VSS inv
    Xi6 IN<6> OUT<6> VDD VSS inv
    Xi5 IN<5> OUT<5> VDD VSS inv
    Xi4 IN<4> OUT<4> VDD VSS inv
    Xi3 IN<3> OUT<3> VDD VSS inv
    Xi2 IN<2> OUT<2> VDD VSS inv
    Xi1 IN<1> OUT<1> VDD VSS inv
    Xi0 IN<0> OUT<0> VDD VSS inv
.ENDS

.SUBCKT cal_tdc_v0 CAL_ENABLE CONF<0> CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> OUT0
                   + OUT1 OUT2 RO_ENABLE RO_OUT RST RST' SEL<0> SEL<1> VDD VSS
    Xi0 net6<0> net6<1> net6<2> net6<3> net6<4> net6<5> net6<6> net6<7> CONF<0> CONF<1> CONF<2>
        + CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> RO_ENABLE RO<0> VDD VSS ro_2i
    Xi1 RO<0> RO<1> RO<2> RO<3> RST RST' VDD VSS freqscaler3
    Xi8 net023 OUT0_I VDD VSS inv_sd
    Xi4 RO<0> RO<1> RO<2> RO<3> MUX_OUT SEL<0> SEL<1> VDD VSS mux4
    Xi5 CONF<0> CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> net6<0> net6<1> net6<2>
        + net6<3> net6<4> net6<5> net6<6> net6<7> VDD VSS inv_bank_8
    Xi7 CAL_ENABLE net027 net023 RST RST' VDD VSS dff_st_ar_dh
    Xi3 RO_OUT OUT1_I OUT2_I net11 RST RST' VDD VSS dff_st_ar_buf
    Xi2 RO_OUT CAL_ENABLE OUT1_I net17 RST RST' VDD VSS dff_st_ar_buf
    Xi12 OUT2_I OUT2 VDD VSS buffer
    Xi11 OUT1_I OUT1 VDD VSS buffer
    Xi10 OUT0_I OUT0 VDD VSS buffer
    Xi9 MUX_OUT RO_OUT VDD VSS buffer
.ENDS

.SUBCKT synchronizer CLK IN OUT RST RST' VDD VSS
    Xi1 CLK net18 OUT net16 RST RST' VDD VSS dff_st_ar_buf
    Xi0 CLK IN net18 net19 RST RST' VDD VSS dff_st_ar_buf
.ENDS

.SUBCKT equalto52 EQUAL IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> VDD VSS
    Xi4 IN<0> IN'<0> VDD VSS inv
    Xi3 IN<1> IN'<1> VDD VSS inv
    Xi2 IN<3> IN'<3> VDD VSS inv
    Xi1 IN<6> IN'<6> VDD VSS inv
    Xi0 IN<7> IN'<7> VDD VSS inv
    Xi6 IN'<3> IN<2> IN'<1> IN'<0> net7 VDD VSS nand4
    Xi5 IN'<7> IN'<6> IN<5> IN<4> net8 VDD VSS nand4
    Xi7 net8 net7 EQUAL VDD VSS nor2
.ENDS

.SUBCKT xnor2 IN0 IN1 OUT VDD VSS
    Mm3 OUT IN0' net20 VDD p_mos l=60n w=240.0n m=1
    Mm2 net20 IN1' VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN0 net21 VDD p_mos l=60n w=240.0n m=1
    Mm0 net21 IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm7 net19 IN1' VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 net18 IN1 VSS VSS n_mos l=60n w=120.0n m=1
    Mm5 OUT IN0' net18 VSS n_mos l=60n w=120.0n m=1
    Mm4 OUT IN0 net19 VSS n_mos l=60n w=120.0n m=1
    Xi1 IN1 IN1' VDD VSS inv
    Xi0 IN0 IN0' VDD VSS inv
.ENDS

.SUBCKT checkequal_8 EQUAL IN0<0> IN0<1> IN0<2> IN0<3> IN0<4> IN0<5> IN0<6> IN0<7> IN1<0> IN1<1>
                     + IN1<2> IN1<3> IN1<4> IN1<5> IN1<6> IN1<7> VDD VSS
    Xi9 IN0<4> IN1<4> XNOR<4> VDD VSS xnor2
    Xi7 IN0<7> IN1<7> XNOR<7> VDD VSS xnor2
    Xi6 IN0<6> IN1<6> XNOR<6> VDD VSS xnor2
    Xi5 IN0<5> IN1<5> XNOR<5> VDD VSS xnor2
    Xi3 IN0<3> IN1<3> XNOR<3> VDD VSS xnor2
    Xi2 IN0<2> IN1<2> XNOR<2> VDD VSS xnor2
    Xi1 IN0<1> IN1<1> XNOR<1> VDD VSS xnor2
    Xi0 IN0<0> IN1<0> XNOR<0> VDD VSS xnor2
    Xi8 XNOR<4> XNOR<5> XNOR<6> XNOR<7> NAND1 VDD VSS nand4
    Xi4 XNOR<0> XNOR<1> XNOR<2> XNOR<3> NAND0 VDD VSS nand4
    Xi10 NAND0 NAND1 EQUAL VDD VSS nor2
.ENDS

.SUBCKT checkequal_16 EQUAL IN0<0> IN0<1> IN0<2> IN0<3> IN0<4> IN0<5> IN0<6> IN0<7> IN0<8> IN0<9>
                      + IN0<10> IN0<11> IN0<12> IN0<13> IN0<14> IN0<15> IN1<0> IN1<1> IN1<2> IN1<3>
                      + IN1<4> IN1<5> IN1<6> IN1<7> IN1<8> IN1<9> IN1<10> IN1<11> IN1<12> IN1<13>
                      + IN1<14> IN1<15> VDD VSS
    Xi1 EQ1 IN0<8> IN0<9> IN0<10> IN0<11> IN0<12> IN0<13> IN0<14> IN0<15> IN1<8> IN1<9> IN1<10>
        + IN1<11> IN1<12> IN1<13> IN1<14> IN1<15> VDD VSS checkequal_8
    Xi0 EQ0 IN0<0> IN0<1> IN0<2> IN0<3> IN0<4> IN0<5> IN0<6> IN0<7> IN1<0> IN1<1> IN1<2> IN1<3>
        + IN1<4> IN1<5> IN1<6> IN1<7> VDD VSS checkequal_8
    Xi2 EQ0 EQ1 net3 VDD VSS nand2
    Xi3 net3 EQUAL VDD VSS inv
.ENDS

.SUBCKT shiftreg_4 CLK IN<0> IN<1> IN<2> IN<3> IN_SER OUT RST RST' SEL_SER VDD VSS
    Xi7 IN<0> IN_SER net3 SEL_SER VDD VSS mux2
    Xi6 IN<1> INT<0> net42 SEL_SER VDD VSS mux2
    Xi5 IN<2> INT<1> net35 SEL_SER VDD VSS mux2
    Xi4 IN<3> INT<2> net17 SEL_SER VDD VSS mux2
    Xi9 CLK net42 INT<1> net40 RST RST' VDD VSS dff_st_ar
    Xi10 CLK net35 INT<2> net32 RST RST' VDD VSS dff_st_ar
    Xi11 CLK net17 OUT net24 RST RST' VDD VSS dff_st_ar
    Xi8 CLK net3 INT<0> net45 RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT shiftreg_8 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN_SER OUT RST RST' SEL_SER
                   + VDD VSS
    Xi1 CLK IN<4> IN<5> IN<6> IN<7> net3 OUT RST RST' SEL_SER VDD VSS shiftreg_4
    Xi0 CLK IN<0> IN<1> IN<2> IN<3> IN_SER net3 RST RST' SEL_SER VDD VSS shiftreg_4
.ENDS

.SUBCKT shiftreg_16 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11>
                    + IN<12> IN<13> IN<14> IN<15> IN_SER OUT RST RST' SEL_SER VDD VSS
    Xi1 CLK IN<8> IN<9> IN<10> IN<11> IN<12> IN<13> IN<14> IN<15> net016 OUT RST RST' SEL_SER VDD
        + VSS shiftreg_8
    Xi0 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN_SER net016 RST RST' SEL_SER VDD VSS
        + shiftreg_8
.ENDS

.SUBCKT shiftreg_52 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11>
                    + IN<12> IN<13> IN<14> IN<15> IN<16> IN<17> IN<18> IN<19> IN<20> IN<21> IN<22>
                    + IN<23> IN<24> IN<25> IN<26> IN<27> IN<28> IN<29> IN<30> IN<31> IN<32> IN<33>
                    + IN<34> IN<35> IN<36> IN<37> IN<38> IN<39> IN<40> IN<41> IN<42> IN<43> IN<44>
                    + IN<45> IN<46> IN<47> IN<48> IN<49> IN<50> IN<51> IN_SER OUT RST RST' SEL_SER
                    + VDD VSS
    Xi2 CLK IN<32> IN<33> IN<34> IN<35> IN<36> IN<37> IN<38> IN<39> IN<40> IN<41> IN<42> IN<43>
        + IN<44> IN<45> IN<46> IN<47> net6 net7 RST RST' SEL_SER VDD VSS shiftreg_16
    Xi1 CLK IN<16> IN<17> IN<18> IN<19> IN<20> IN<21> IN<22> IN<23> IN<24> IN<25> IN<26> IN<27>
        + IN<28> IN<29> IN<30> IN<31> net5 net6 RST RST' SEL_SER VDD VSS shiftreg_16
    Xi0 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11> IN<12> IN<13>
        + IN<14> IN<15> IN_SER net5 RST RST' SEL_SER VDD VSS shiftreg_16
    Xi3 CLK IN<48> IN<49> IN<50> IN<51> net7 OUT RST RST' SEL_SER VDD VSS shiftreg_4
.ENDS

.SUBCKT conf_datapath CAL_EN CAL_OUT0 CAL_OUT1 CAL_OUT2 CAL_ROOUT CAL_RO_EN CLK CONF_STATECNT<0>
                      + CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4>
                      + CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8>
                      + CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12>
                      + CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> CONF_TDCCAL<0>
                      + CONF_TDCCAL<1> CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4> CONF_TDCCAL<5>
                      + CONF_TDCCAL<6> CONF_TDCCAL<7> CONF_TDCCAL<8> CONF_TDCCAL<9> DATA_OUT
                      + DATA_READY RST RST' SEND_DATA<32> SEND_DATA<33> SEND_DATA<34> SEND_DATA<35>
                      + SEND_DATA<36> SEND_DATA<37> SEND_DATA<38> SEND_DATA<39> SEND_DATA<40>
                      + SEND_DATA<41> SEND_DATA<42> SEND_DATA<43> SEND_DATA<44> SEND_DATA<45>
                      + SEND_DATA<46> SEND_DATA<47> SEND_DATA<48> SEND_DATA<49> SEND_DATA<50>
                      + SEND_DATA<51> SER_CLK SER_READY STA_READY TDC0_INT TDC0_READY TDC1_INT
                      + TDC1_READY TDC_READY VDD VSS
    Xi3 CLK STATE_CNT<0> STATE_CNT<1> STATE_CNT<2> STATE_CNT<3> STATE_CNT<4> STATE_CNT<5>
        + STATE_CNT<6> STATE_CNT<7> STATE_CNT<8> STATE_CNT<9> STATE_CNT<10> STATE_CNT<11>
        + STATE_CNT<12> STATE_CNT<13> STATE_CNT<14> STATE_CNT<15> net010 RST RST' VDD VSS
        + asynccounter_16
    Xi1 TDC0_INT SEND_DATA<0> SEND_DATA<1> SEND_DATA<2> SEND_DATA<3> SEND_DATA<4> SEND_DATA<5>
        + SEND_DATA<6> SEND_DATA<7> SEND_DATA<8> SEND_DATA<9> SEND_DATA<10> SEND_DATA<11>
        + SEND_DATA<12> SEND_DATA<13> SEND_DATA<14> SEND_DATA<15> net7 RST RST' VDD VSS
        + asynccounter_16
    Xi0 TDC1_INT SEND_DATA<16> SEND_DATA<17> SEND_DATA<18> SEND_DATA<19> SEND_DATA<20> SEND_DATA<21>
        + SEND_DATA<22> SEND_DATA<23> SEND_DATA<24> SEND_DATA<25> SEND_DATA<26> SEND_DATA<27>
        + SEND_DATA<28> SEND_DATA<29> SEND_DATA<30> SEND_DATA<31> net10 RST RST' VDD VSS
        + asynccounter_16
    Xi2 CAL_EN CONF_TDCCAL<0> CONF_TDCCAL<1> CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4>
        + CONF_TDCCAL<5> CONF_TDCCAL<6> CONF_TDCCAL<7> CAL_OUT0 CAL_OUT1 CAL_OUT2 CAL_RO_EN
        + CAL_ROOUT RST RST' CONF_TDCCAL<8> CONF_TDCCAL<9> VDD VSS cal_tdc_v0
    Xi4 net03 SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> net028 RST RST' VDD VSS asynccounter_8
    Xi10 CLK TDC0_READY TDC0_READYSYNC RST RST' VDD VSS synchronizer
    Xi9 CLK TDC1_READY TDC1_READYSYNC RST RST' VDD VSS synchronizer
    Xi5 CLK SER_CLK net03 RST RST' VDD VSS synchronizer
    Xi7 SER_READY SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> VDD VSS equalto52
    Xi8 STA_READY STATE_CNT<0> STATE_CNT<1> STATE_CNT<2> STATE_CNT<3> STATE_CNT<4> STATE_CNT<5>
        + STATE_CNT<6> STATE_CNT<7> STATE_CNT<8> STATE_CNT<9> STATE_CNT<10> STATE_CNT<11>
        + STATE_CNT<12> STATE_CNT<13> STATE_CNT<14> STATE_CNT<15> CONF_STATECNT<0> CONF_STATECNT<1>
        + CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6>
        + CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11>
        + CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> VDD VSS
        + checkequal_16
    Xi11 TDC0_READYSYNC TDC1_READYSYNC net09 VDD VSS nand2
    Xi12 net09 TDC_READY VDD VSS inv
    Xi13 Shift_CLK SEND_DATA<0> SEND_DATA<1> SEND_DATA<2> SEND_DATA<3> SEND_DATA<4> SEND_DATA<5>
         + SEND_DATA<6> SEND_DATA<7> SEND_DATA<8> SEND_DATA<9> SEND_DATA<10> SEND_DATA<11>
         + SEND_DATA<12> SEND_DATA<13> SEND_DATA<14> SEND_DATA<15> SEND_DATA<16> SEND_DATA<17>
         + SEND_DATA<18> SEND_DATA<19> SEND_DATA<20> SEND_DATA<21> SEND_DATA<22> SEND_DATA<23>
         + SEND_DATA<24> SEND_DATA<25> SEND_DATA<26> SEND_DATA<27> SEND_DATA<28> SEND_DATA<29>
         + SEND_DATA<30> SEND_DATA<31> SEND_DATA<32> SEND_DATA<33> SEND_DATA<34> SEND_DATA<35>
         + SEND_DATA<36> SEND_DATA<37> SEND_DATA<38> SEND_DATA<39> SEND_DATA<40> SEND_DATA<41>
         + SEND_DATA<42> SEND_DATA<43> SEND_DATA<44> SEND_DATA<45> SEND_DATA<46> SEND_DATA<47>
         + SEND_DATA<48> SEND_DATA<49> SEND_DATA<50> SEND_DATA<51> SEND_DATA<0> DATA_OUT RST RST'
         + DATA_READY VDD VSS shiftreg_52
    Xi14 CLK SER_CLK Shift_CLK DATA_READY VDD VSS mux2
.ENDS

.SUBCKT conf_toplevel CAL_EN CAL_OUT0 CAL_OUT1 CAL_OUT2 CAL_ROOUT CAL_RO_EN CLK CONF_STATECNT<0>
                      + CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4>
                      + CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8>
                      + CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12>
                      + CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> CONF_TDCCAL<0>
                      + CONF_TDCCAL<1> CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4> CONF_TDCCAL<5>
                      + CONF_TDCCAL<6> CONF_TDCCAL<7> CONF_TDCCAL<8> CONF_TDCCAL<9> DATA_OUT
                      + DATA_READY DAT_RST DAT_RST' RST RST' SER_CLK SER_READY STATE<0> STATE<1>
                      + STATE<2> STA_READY TDC0_ALARM<0> TDC0_ALARM<1> TDC0_FF<0> TDC0_FF<1>
                      + TDC0_FF<2> TDC0_FF<3> TDC0_FF<4> TDC0_FF<5> TDC0_FF<6> TDC0_FF<7> TDC0_INT
                      + TDC0_READY TDC1_ALARM<0> TDC1_ALARM<1> TDC1_FF<0> TDC1_FF<1> TDC1_FF<2>
                      + TDC1_FF<3> TDC1_FF<4> TDC1_FF<5> TDC1_FF<6> TDC1_FF<7> TDC1_INT TDC1_READY
                      + TDC_READY VDD VSS
    Xi0 CAL_EN CAL_RO_EN CLK CTRL_RST DATA_READY RST RST' SER_READY STATE<0> STATE<1> STATE<2>
        + STA_READY TDC_READY VDD VSS conf_control
    Xi1 CAL_EN CAL_OUT0 CAL_OUT1 CAL_OUT2 CAL_ROOUT CAL_RO_EN CLK CONF_STATECNT<0> CONF_STATECNT<1>
        + CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6>
        + CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11>
        + CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> CONF_TDCCAL<0>
        + CONF_TDCCAL<1> CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4> CONF_TDCCAL<5> CONF_TDCCAL<6>
        + CONF_TDCCAL<7> CONF_TDCCAL<8> CONF_TDCCAL<9> DATA_OUT DATA_READY DAT_RST DAT_RST'
        + TDC0_FF<0> TDC0_FF<1> TDC0_FF<2> TDC0_FF<3> TDC0_FF<4> TDC0_FF<5> TDC0_FF<6> TDC0_FF<7>
        + TDC1_FF<0> TDC1_FF<1> TDC1_FF<2> TDC1_FF<3> TDC1_FF<4> TDC1_FF<5> TDC1_FF<6> TDC1_FF<7>
        + TDC0_ALARM<0> TDC0_ALARM<1> TDC1_ALARM<0> TDC1_ALARM<1> SER_CLK SER_READY STA_READY
        + TDC0_INT TDC0_READY TDC1_INT TDC1_READY TDC_READY VDD VSS conf_datapath
    Xi2 CTRL_RST CTRL_RST' VDD VSS inv
    Xi3 CTRL_RST RST DAT_RST_INT' VDD VSS nor2
    Xi4 CTRL_RST' RST' DAT_RST_INT VDD VSS nand2
    Xi6 DAT_RST_INT DAT_RST VDD VSS buffer
    Xi5 DAT_RST_INT' DAT_RST' VDD VSS buffer
.ENDS

.SUBCKT equalto24 EQUAL IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> VDD VSS
    Xi5 IN<7> IN'<7> VDD VSS inv
    Xi4 IN<6> IN'<6> VDD VSS inv
    Xi3 IN<5> IN'<5> VDD VSS inv
    Xi2 IN<2> IN'<2> VDD VSS inv
    Xi1 IN<1> IN'<1> VDD VSS inv
    Xi0 IN<0> IN'<0> VDD VSS inv
    Xi7 IN<4> IN'<5> IN'<6> IN'<7> net11 VDD VSS nand4
    Xi6 IN'<0> IN'<1> IN'<2> IN<3> net12 VDD VSS nand4
    Xi8 net12 net11 EQUAL VDD VSS nor2
.ENDS

.SUBCKT shiftreg_24 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11>
                    + IN<12> IN<13> IN<14> IN<15> IN<16> IN<17> IN<18> IN<19> IN<20> IN<21> IN<22>
                    + IN<23> IN_SER OUT RST RST' SEL_SER VDD VSS
    Xi0 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN_SER net17 RST RST' SEL_SER VDD VSS
        + shiftreg_8
    Xi1 CLK IN<8> IN<9> IN<10> IN<11> IN<12> IN<13> IN<14> IN<15> IN<16> IN<17> IN<18> IN<19> IN<20>
        + IN<21> IN<22> IN<23> net17 OUT RST RST' SEL_SER VDD VSS shiftreg_16
.ENDS

.SUBCKT bit_datapath CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3>
                     + CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7>
                     + CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11>
                     + CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15>
                     + DATA_OUT DATA_READY DC_INT RST RST' SEND_DATA<0> SEND_DATA<1> SEND_DATA<2>
                     + SEND_DATA<3> SEND_DATA<4> SEND_DATA<5> SEND_DATA<6> SEND_DATA<7> SER_CLK
                     + SER_READY STA_READY TDC0_READY TDC1_READY TDC_READY VDD VSS
    Xi10 CLK STA_CNT<0> STA_CNT<1> STA_CNT<2> STA_CNT<3> STA_CNT<4> STA_CNT<5> STA_CNT<6> STA_CNT<7>
         + STA_CNT<8> STA_CNT<9> STA_CNT<10> STA_CNT<11> STA_CNT<12> STA_CNT<13> STA_CNT<14>
         + STA_CNT<15> net030 RST RST' VDD VSS asynccounter_16
    Xi0 DC_INT SEND_DATA<8> SEND_DATA<9> SEND_DATA<10> SEND_DATA<11> SEND_DATA<12> SEND_DATA<13>
        + SEND_DATA<14> SEND_DATA<15> SEND_DATA<16> SEND_DATA<17> SEND_DATA<18> SEND_DATA<19>
        + SEND_DATA<20> SEND_DATA<21> SEND_DATA<22> SEND_DATA<23> net7 RST RST' VDD VSS
        + asynccounter_16
    Xi6 CLK TDC1_READY TDC1_READY_S RST RST' VDD VSS synchronizer
    Xi5 CLK TDC0_READY TDC0_READY_S RST RST' VDD VSS synchronizer
    Xi1 CLK SER_CLK net10 RST RST' VDD VSS synchronizer
    Xi2 net10 SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> net15 RST RST' VDD VSS asynccounter_8
    Xi3 SER_READY SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> VDD VSS equalto24
    Xi4 Shift_CLK SEND_DATA<0> SEND_DATA<1> SEND_DATA<2> SEND_DATA<3> SEND_DATA<4> SEND_DATA<5>
        + SEND_DATA<6> SEND_DATA<7> SEND_DATA<8> SEND_DATA<9> SEND_DATA<10> SEND_DATA<11>
        + SEND_DATA<12> SEND_DATA<13> SEND_DATA<14> SEND_DATA<15> SEND_DATA<16> SEND_DATA<17>
        + SEND_DATA<18> SEND_DATA<19> SEND_DATA<20> SEND_DATA<21> SEND_DATA<22> SEND_DATA<23>
        + SEND_DATA<0> DATA_OUT RST RST' DATA_READY VDD VSS shiftreg_24
    Xi7 TDC0_READY_S TDC1_READY_S net038 VDD VSS nand2
    Xi8 net038 TDC_READY VDD VSS inv
    Xi9 CLK SER_CLK Shift_CLK DATA_READY VDD VSS mux2
    Xi11 STA_READY STA_CNT<0> STA_CNT<1> STA_CNT<2> STA_CNT<3> STA_CNT<4> STA_CNT<5> STA_CNT<6>
         + STA_CNT<7> STA_CNT<8> STA_CNT<9> STA_CNT<10> STA_CNT<11> STA_CNT<12> STA_CNT<13>
         + STA_CNT<14> STA_CNT<15> CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2>
         + CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7>
         + CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12>
         + CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> VDD VSS checkequal_16
.ENDS

.SUBCKT bit_toplevel ALARM_DC CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2>
                     + CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6>
                     + CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10>
                     + CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
                     + CONF_STATECNT<15> DATA_OUT DATA_READY DAT_RST DAT_RST' DC_INT E2L_EN MERO_EN
                     + RAND0 RAND1 RST RST' SEND_FREE SER_CLK SER_READY STATE<0> STATE<1> STATE<2>
                     + STA_READY TDC0_ALARM<0> TDC0_ALARM<1> TDC0_READY TDC1_ALARM<0> TDC1_ALARM<1>
                     + TDC1_READY TDC_READY VDD VSS
    Xi0 CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4>
        + CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9>
        + CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
        + CONF_STATECNT<15> DATA_OUT DATA_READY DC_INT DAT_RST DAT_RST' TDC0_ALARM<0> TDC0_ALARM<1>
        + TDC1_ALARM<0> TDC1_ALARM<1> ALARM_DC RAND0 RAND1 SEND_FREE SER_CLK SER_READY STA_READY
        + TDC0_READY TDC1_READY TDC_READY VDD VSS bit_datapath
    Xi1 E2L_EN MERO_EN CLK CTRL_RST DATA_READY RST RST' SER_READY STATE<0> STATE<1> STATE<2>
        + STA_READY TDC_READY VDD VSS conf_control
    Xi2 CTRL_RST CTRL_RST' VDD VSS inv
    Xi3 CTRL_RST' RST' DAT_RST_I VDD VSS nand2
    Xi4 CTRL_RST RST DAT_RST_I' VDD VSS nor2
    Xi6 DAT_RST_I' DAT_RST' VDD VSS buffer
    Xi5 DAT_RST_I DAT_RST VDD VSS buffer
.ENDS

.SUBCKT async_control_0 CLK MERO_E2L MERO_EN RST RST' STATE<0> STATE<1> STA_READY TDC_READY TRNG_RST
                        + VDD VSS
    Xi1 CLK NEXTSTATE<1> STATE<1> TRNG_RST RST RST' VDD VSS dff_st_ar
    Xi0 CLK NEXTSTATE<0> STATE<0> STATE'<0> RST RST' VDD VSS dff_st_ar
    Xi8 STATE'<0> STATE<1> net08 VDD VSS nand2
    Xi7 STATE1_INT STATE'<0> NEXTSTATE<1> VDD VSS nand2
    Xi6 STATE<1> TDC_READY' STATE1_INT VDD VSS nand2
    Xi3 STATE0_INT STATE<1> NEXTSTATE<0> VDD VSS nand2
    Xi2 STATE<0> STA_READY' STATE0_INT VDD VSS nand2
    Xi9 net08 MERO_E2L_I VDD VSS inv
    Xi5 TDC_READY TDC_READY' VDD VSS inv
    Xi4 STA_READY STA_READY' VDD VSS inv
    Xi11 STATE<1> MERO_EN VDD VSS buffer
    Xi10 MERO_E2L_I MERO_E2L VDD VSS buffer
.ENDS

.SUBCKT async_control_1 CLK CLK_EN CLK_READY CTRL_RST DATA_READY RST RST' SER_READY STATE<0>
                        + STATE<1> STATE<2> VDD VSS
    Xi2 CLK NEXTSTATE<2> STATE<2> STATE'<2> RST RST' VDD VSS dff_st_ar
    Xi1 CLK NEXTSTATE<1> STATE<1> STATE'<1> RST RST' VDD VSS dff_st_ar
    Xi0 CLK NEXTSTATE<0> STATE<0> STATE'<0> RST RST' VDD VSS dff_st_ar
    Xi15 STATE'<1> STATE'<2> DATA_READY_I VDD VSS nor2
    Xi13 STATE<1> STATE<2> CLK_EN_I VDD VSS nor2
    Xi3 STATE<1> STATE<2> NEXTSTATE<0> VDD VSS nor2
    Xi9 STATE'<0> STATE<1> net05 VDD VSS nand2
    Xi7 STATE<0> CLK_READY STATE1_INT<3> VDD VSS nand2
    Xi6 STATE<1> STATE'<2> STATE1_INT<2> VDD VSS nand2
    Xi5 STATE<0> STATE<1> STATE1_INT<1> VDD VSS nand2
    Xi4 STATE<1> SER_READY' STATE1_INT<0> VDD VSS nand2
    Xi8 STATE1_INT<0> STATE1_INT<1> STATE1_INT<2> STATE1_INT<3> NEXTSTATE<1> VDD VSS nand4
    Xi11 SER_READY SER_READY' VDD VSS inv
    Xi10 net05 NEXTSTATE<2> VDD VSS inv
    Xi14 STATE<0> STATE<1> STATE<2> CTRL_RST VDD VSS nor3
    Xi17 DATA_READY_I DATA_READY VDD VSS buffer
    Xi16 CLK_EN_I CLK_EN VDD VSS buffer
.ENDS

.SUBCKT asynccounterequal_16 CLK CONF_EQUAL<0> CONF_EQUAL<1> CONF_EQUAL<2> CONF_EQUAL<3>
                             + CONF_EQUAL<4> CONF_EQUAL<5> CONF_EQUAL<6> CONF_EQUAL<7> CONF_EQUAL<8>
                             + CONF_EQUAL<9> CONF_EQUAL<10> CONF_EQUAL<11> CONF_EQUAL<12>
                             + CONF_EQUAL<13> CONF_EQUAL<14> CONF_EQUAL<15> EQUAL RST RST' VDD VSS
    Xi0 CLK CNT<0> CNT<1> CNT<2> CNT<3> CNT<4> CNT<5> CNT<6> CNT<7> CNT<8> CNT<9> CNT<10> CNT<11>
        + CNT<12> CNT<13> CNT<14> CNT<15> net13 RST RST' VDD VSS asynccounter_16
    Xi1 EQUAL CNT<0> CNT<1> CNT<2> CNT<3> CNT<4> CNT<5> CNT<6> CNT<7> CNT<8> CNT<9> CNT<10> CNT<11>
        + CNT<12> CNT<13> CNT<14> CNT<15> CONF_EQUAL<0> CONF_EQUAL<1> CONF_EQUAL<2> CONF_EQUAL<3>
        + CONF_EQUAL<4> CONF_EQUAL<5> CONF_EQUAL<6> CONF_EQUAL<7> CONF_EQUAL<8> CONF_EQUAL<9>
        + CONF_EQUAL<10> CONF_EQUAL<11> CONF_EQUAL<12> CONF_EQUAL<13> CONF_EQUAL<14> CONF_EQUAL<15>
        + VDD VSS checkequal_16
.ENDS

.SUBCKT async_datapath_0 CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3>
                         + CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7>
                         + CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11>
                         + CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15>
                         + RST RST' STA_READY TDC0_READY TDC1_READY TDC_READY VDD VSS
    Xi1 CLK TDC1_READY TDC1_SYNC RST RST' VDD VSS synchronizer
    Xi0 CLK TDC0_READY TDC0_SYNC RST RST' VDD VSS synchronizer
    Xi2 TDC0_SYNC TDC1_SYNC net7 VDD VSS nand2
    Xi3 net7 TDC_READY VDD VSS inv
    Xi5 CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4>
        + CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9>
        + CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
        + CONF_STATECNT<15> STA_READY RST RST' VDD VSS asynccounterequal_16
.ENDS

.SUBCKT asynccounter_32 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                        + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18>
                        + OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27>
                        + OUT<28> OUT<29> OUT<30> OUT<31> Q' RST RST' VDD VSS
    Xi1 net7 OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26>
        + OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> Q' RST RST' VDD VSS asynccounter_16
    Xi0 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10> OUT<11>
        + OUT<12> OUT<13> OUT<14> OUT<15> net7 RST RST' VDD VSS asynccounter_16
.ENDS

.SUBCKT shiftreg_32 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11>
                    + IN<12> IN<13> IN<14> IN<15> IN<16> IN<17> IN<18> IN<19> IN<20> IN<21> IN<22>
                    + IN<23> IN<24> IN<25> IN<26> IN<27> IN<28> IN<29> IN<30> IN<31> IN_SER OUT RST
                    + RST' SEL_SER VDD VSS
    Xi1 CLK IN<16> IN<17> IN<18> IN<19> IN<20> IN<21> IN<22> IN<23> IN<24> IN<25> IN<26> IN<27>
        + IN<28> IN<29> IN<30> IN<31> net7 OUT RST RST' SEL_SER VDD VSS shiftreg_16
    Xi0 CLK IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11> IN<12> IN<13>
        + IN<14> IN<15> IN_SER net7 RST RST' SEL_SER VDD VSS shiftreg_16
.ENDS

.SUBCKT equalto32 EQUAL IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> VDD VSS
    Xi8 IN<4> IN'<4> VDD VSS inv
    Xi7 IN<6> IN'<6> VDD VSS inv
    Xi6 IN<7> IN'<7> VDD VSS inv
    Xi5 IN<3> IN'<3> VDD VSS inv
    Xi3 IN<1> IN'<1> VDD VSS inv
    Xi4 IN<2> IN'<2> VDD VSS inv
    Xi0 IN<0> IN'<0> VDD VSS inv
    Xi10 IN'<4> IN<5> IN'<6> IN'<7> net013 VDD VSS nand4
    Xi9 IN'<0> IN'<1> IN'<2> IN'<3> net014 VDD VSS nand4
    Xi11 net014 net013 EQUAL VDD VSS nor2
.ENDS

.SUBCKT async_datapath_1 CLK CLK_EN CLK_READY CONF_TDCCNT<0> CONF_TDCCNT<1> CONF_TDCCNT<2>
                         + CONF_TDCCNT<3> CONF_TDCCNT<4> CONF_TDCCNT<5> CONF_TDCCNT<6>
                         + CONF_TDCCNT<7> CONF_TDCCNT<8> CONF_TDCCNT<9> CONF_TDCCNT<10>
                         + CONF_TDCCNT<11> CONF_TDCCNT<12> CONF_TDCCNT<13> CONF_TDCCNT<14>
                         + CONF_TDCCNT<15> DATA_OUT DATA_READY RST RST' SER_CLK SER_READY TDC_READY
                         + VDD VSS
    Xi0 TDC_READY CONF_TDCCNT<0> CONF_TDCCNT<1> CONF_TDCCNT<2> CONF_TDCCNT<3> CONF_TDCCNT<4>
        + CONF_TDCCNT<5> CONF_TDCCNT<6> CONF_TDCCNT<7> CONF_TDCCNT<8> CONF_TDCCNT<9> CONF_TDCCNT<10>
        + CONF_TDCCNT<11> CONF_TDCCNT<12> CONF_TDCCNT<13> CONF_TDCCNT<14> CONF_TDCCNT<15> CLK_READY
        + RST RST' VDD VSS asynccounterequal_16
    Xi1 net04 CLK_CNT<0> CLK_CNT<1> CLK_CNT<2> CLK_CNT<3> CLK_CNT<4> CLK_CNT<5> CLK_CNT<6>
        + CLK_CNT<7> CLK_CNT<8> CLK_CNT<9> CLK_CNT<10> CLK_CNT<11> CLK_CNT<12> CLK_CNT<13>
        + CLK_CNT<14> CLK_CNT<15> CLK_CNT<16> CLK_CNT<17> CLK_CNT<18> CLK_CNT<19> CLK_CNT<20>
        + CLK_CNT<21> CLK_CNT<22> CLK_CNT<23> CLK_CNT<24> CLK_CNT<25> CLK_CNT<26> CLK_CNT<27>
        + CLK_CNT<28> CLK_CNT<29> CLK_CNT<30> CLK_CNT<31> net09 RST RST' VDD VSS asynccounter_32
    Xi2 CLK CLK_EN net05 VDD VSS nand2
    Xi3 net05 net04 VDD VSS inv
    Xi4 SHIFT_CLK CLK_CNT<0> CLK_CNT<1> CLK_CNT<2> CLK_CNT<3> CLK_CNT<4> CLK_CNT<5> CLK_CNT<6>
        + CLK_CNT<7> CLK_CNT<8> CLK_CNT<9> CLK_CNT<10> CLK_CNT<11> CLK_CNT<12> CLK_CNT<13>
        + CLK_CNT<14> CLK_CNT<15> CLK_CNT<16> CLK_CNT<17> CLK_CNT<18> CLK_CNT<19> CLK_CNT<20>
        + CLK_CNT<21> CLK_CNT<22> CLK_CNT<23> CLK_CNT<24> CLK_CNT<25> CLK_CNT<26> CLK_CNT<27>
        + CLK_CNT<28> CLK_CNT<29> CLK_CNT<30> CLK_CNT<31> CLK_CNT<0> DATA_OUT RST RST' DATA_READY
        + VDD VSS shiftreg_32
    Xi5 CLK SER_CLK net021 DATA_READY VDD VSS mux2
    Xi6 CLK SER_CLK net027 RST RST' VDD VSS synchronizer
    Xi7 net027 SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> net025 RST RST' VDD VSS asynccounter_8
    Xi8 SER_READY SER_CNT<0> SER_CNT<1> SER_CNT<2> SER_CNT<3> SER_CNT<4> SER_CNT<5> SER_CNT<6>
        + SER_CNT<7> VDD VSS equalto32
    Xi9 net021 SHIFT_CLK VDD VSS buffer
.ENDS

.SUBCKT async_toplevel CLK CLK_EN CLK_READY CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2>
                       + CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6>
                       + CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10>
                       + CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
                       + CONF_STATECNT<15> CONF_TDCCNT<0> CONF_TDCCNT<1> CONF_TDCCNT<2>
                       + CONF_TDCCNT<3> CONF_TDCCNT<4> CONF_TDCCNT<5> CONF_TDCCNT<6> CONF_TDCCNT<7>
                       + CONF_TDCCNT<8> CONF_TDCCNT<9> CONF_TDCCNT<10> CONF_TDCCNT<11>
                       + CONF_TDCCNT<12> CONF_TDCCNT<13> CONF_TDCCNT<14> CONF_TDCCNT<15> DATA_OUT
                       + DATA_READY DP0_RST DP0_RST' DP1_RST MERO_E2L MERO_EN RST RST' SER_CLK
                       + SER_READY STATE0<0> STATE0<1> STATE1<0> STATE1<1> STATE1<2> STA_READY
                       + TDC0_READY TDC1_READY TDC_READY VDD VSS
    Xi0 CLK MERO_E2L MERO_EN RST RST' STATE0<0> STATE0<1> STA_READY TDC_READY CTRL0_RST VDD VSS
        + async_control_0
    Xi1 CLK CLK_EN CLK_READY CTRL1_RST DATA_READY RST RST' SER_READY STATE1<0> STATE1<1> STATE1<2>
        + VDD VSS async_control_1
    Xi2 CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4>
        + CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9>
        + CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
        + CONF_STATECNT<15> DP0_RST DP0_RST' STA_READY TDC0_READY TDC1_READY TDC_READY VDD VSS
        + async_datapath_0
    Xi3 CLK CLK_EN CLK_READY CONF_TDCCNT<0> CONF_TDCCNT<1> CONF_TDCCNT<2> CONF_TDCCNT<3>
        + CONF_TDCCNT<4> CONF_TDCCNT<5> CONF_TDCCNT<6> CONF_TDCCNT<7> CONF_TDCCNT<8> CONF_TDCCNT<9>
        + CONF_TDCCNT<10> CONF_TDCCNT<11> CONF_TDCCNT<12> CONF_TDCCNT<13> CONF_TDCCNT<14>
        + CONF_TDCCNT<15> DATA_OUT DATA_READY DP1_RST DP1_RST' SER_CLK SER_READY TDC_READY VDD VSS
        + async_datapath_1
    Xi5 CTRL1_RST' RST' DP1_RST_I VDD VSS nand2
    Xi4 CTRL0_RST' RST' DP0_RST_I VDD VSS nand2
    Xi7 CTRL1_RST RST DP1_RST'_I VDD VSS nor2
    Xi6 CTRL0_RST RST DP0_RST'_I VDD VSS nor2
    Xi11 DP1_RST'_I DP1_RST' VDD VSS buffer
    Xi10 DP1_RST_I DP1_RST VDD VSS buffer
    Xi9 DP0_RST'_I DP0_RST' VDD VSS buffer
    Xi8 DP0_RST_I DP0_RST VDD VSS buffer
    Xi13 CTRL1_RST CTRL1_RST' VDD VSS inv
    Xi12 CTRL0_RST CTRL0_RST' VDD VSS inv
.ENDS

.SUBCKT buffer_large IN OUT VDD VSS
    Mm7 OUT INT<2> VSS VSS n_mos l=60n w=480.0n m=16
    Mm5 INT<2> INT<1> VSS VSS n_mos l=60n w=480.0n m=4
    Mm2 INT<1> INT<0> VSS VSS n_mos l=60n w=480.0n m=1
    Mm0 INT<0> IN VSS VSS n_mos l=60n w=120.0n m=1
    Mm6 OUT INT<2> VDD VDD p_mos l=60n w=480.0n m=16
    Mm4 INT<2> INT<1> VDD VDD p_mos l=60n w=480.0n m=4
    Mm3 INT<1> INT<0> VDD VDD p_mos l=60n w=480.0n m=1
    Mm1 INT<0> IN VDD VDD p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT freq_scaler2 CLK OUT<0> OUT<1> Q' RST RST' VDD VSS
    Xi1 INT OUT<1> Q' RST RST' VDD VSS tff_st_ar
    Xi0 CLK OUT<0> INT RST RST' VDD VSS tff_st_ar
.ENDS

.SUBCKT freq_scaler4 CLK OUT<0> OUT<1> OUT<2> OUT<3> Q' RST RST' VDD VSS
    Xi1 net17 OUT<2> OUT<3> Q' RST RST' VDD VSS freq_scaler2
    Xi0 CLK OUT<0> OUT<1> net17 RST RST' VDD VSS freq_scaler2
.ENDS

.SUBCKT freq_scaler8 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> Q' RST RST' VDD VSS
    Xi1 net17 OUT<4> OUT<5> OUT<6> OUT<7> Q' RST RST' VDD VSS freq_scaler4
    Xi0 CLK OUT<0> OUT<1> OUT<2> OUT<3> net17 RST RST' VDD VSS freq_scaler4
.ENDS

.SUBCKT freq_scaler16 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                      + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> Q' RST RST' VDD VSS
    Xi1 net17 OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> Q' RST RST' VDD VSS
        + freq_scaler8
    Xi0 CLK OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> net17 RST RST' VDD VSS
        + freq_scaler8
.ENDS

.SUBCKT mux16 IN<0> IN<1> IN<2> IN<3> IN<4> IN<5> IN<6> IN<7> IN<8> IN<9> IN<10> IN<11> IN<12>
              + IN<13> IN<14> IN<15> OUT SEL<0> SEL<1> SEL<2> SEL<3> VDD VSS
    Xi4 IN<12> IN<13> IN<14> IN<15> INT<3> SEL<0> SEL<1> VDD VSS mux4
    Xi3 IN<8> IN<9> IN<10> IN<11> INT<2> SEL<0> SEL<1> VDD VSS mux4
    Xi5 INT<0> INT<1> INT<2> INT<3> OUT SEL<2> SEL<3> VDD VSS mux4
    Xi1 IN<4> IN<5> IN<6> IN<7> INT<1> SEL<0> SEL<1> VDD VSS mux4
    Xi0 IN<0> IN<1> IN<2> IN<3> INT<0> SEL<0> SEL<1> VDD VSS mux4
.ENDS

.SUBCKT clkmanager CLK CONF_CLK<0> CONF_CLK<1> CONF_CLK<2> CONF_CLK<3> CONF_CLK<4> CONF_CLK<5>
                   + CONF_CLK<6> CONF_CLK<7> CONF_CLK<8> CONF_CLK<9> CONF_CLK<10> CONF_CLK<11>
                   + ENABLE RST RST' VDD VSS
    Xi0 CONF_CLK'<0> CONF_CLK'<1> CONF_CLK'<2> CONF_CLK'<3> CONF_CLK'<4> CONF_CLK'<5> CONF_CLK'<6>
        + CONF_CLK'<7> CONF_CLK<0> CONF_CLK<1> CONF_CLK<2> CONF_CLK<3> CONF_CLK<4> CONF_CLK<5>
        + CONF_CLK<6> CONF_CLK<7> ENABLE MUX_IN<15> VDD VSS ro_2i
    Xi1 MUX_IN<15> MUX_IN<0> MUX_IN<1> MUX_IN<2> MUX_IN<3> MUX_IN<4> MUX_IN<5> MUX_IN<6> MUX_IN<7>
        + MUX_IN<8> MUX_IN<9> MUX_IN<10> MUX_IN<11> MUX_IN<12> MUX_IN<13> MUX_IN<14> net010 net11
        + RST RST' VDD VSS freq_scaler16
    Xi3 MUX_IN<0> MUX_IN<1> MUX_IN<2> MUX_IN<3> MUX_IN<4> MUX_IN<5> MUX_IN<6> MUX_IN<7> MUX_IN<8>
        + MUX_IN<9> MUX_IN<10> MUX_IN<11> MUX_IN<12> MUX_IN<13> MUX_IN<14> MUX_IN<15> net17
        + CONF_CLK<8> CONF_CLK<9> CONF_CLK<10> CONF_CLK<11> VDD VSS mux16
    Xi2 net17 CLK VDD VSS buffer_large
    Xi4 CONF_CLK<0> CONF_CLK<1> CONF_CLK<2> CONF_CLK<3> CONF_CLK<4> CONF_CLK<5> CONF_CLK<6>
        + CONF_CLK<7> CONF_CLK'<0> CONF_CLK'<1> CONF_CLK'<2> CONF_CLK'<3> CONF_CLK'<4> CONF_CLK'<5>
        + CONF_CLK'<6> CONF_CLK'<7> VDD VSS inv_bank_8
.ENDS

.SUBCKT oneto18 IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
                + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> VDD VSS
    Xi17 IN OUT<9> VDD VSS inv
    Xi16 IN OUT<16> VDD VSS inv
    Xi15 IN OUT<17> VDD VSS inv
    Xi14 IN OUT<15> VDD VSS inv
    Xi13 IN OUT<12> VDD VSS inv
    Xi12 IN OUT<14> VDD VSS inv
    Xi11 IN OUT<13> VDD VSS inv
    Xi10 IN OUT<11> VDD VSS inv
    Xi9 IN OUT<10> VDD VSS inv
    Xi8 IN OUT<7> VDD VSS inv
    Xi7 IN OUT<8> VDD VSS inv
    Xi6 IN OUT<6> VDD VSS inv
    Xi5 IN OUT<3> VDD VSS inv
    Xi4 IN OUT<5> VDD VSS inv
    Xi3 IN OUT<4> VDD VSS inv
    Xi2 IN OUT<2> VDD VSS inv
    Xi1 IN OUT<1> VDD VSS inv
    Xi0 IN OUT<0> VDD VSS inv
.ENDS

.SUBCKT ctrl_trng_combo CONF_CLK<0> CONF_CLK<1> CONF_CLK<2> CONF_CLK<3> CONF_CLK<4> CONF_CLK<5>
                        + CONF_CLK<6> CONF_CLK<7> CONF_CLK<8> CONF_CLK<9> CONF_CLK<10> CONF_CLK<11>
                        + CONF_CLKENABLE CONF_CLKSEL CONF_CTRLSEL<0> CONF_CTRLSEL<1>
                        + CONF_DCEDGESEL<0> CONF_DCEDGESEL<1> CONF_DEC0<0> CONF_DEC0<1> CONF_DEC0<2>
                        + CONF_DEC0<3> CONF_DEC0<4> CONF_DEC0<5> CONF_DEC0<6> CONF_DEC0<7>
                        + CONF_DEC0<8> CONF_DEC0<9> CONF_DEC1<0> CONF_DEC1<1> CONF_DEC1<2>
                        + CONF_DEC1<3> CONF_DEC1<4> CONF_DEC1<5> CONF_DEC1<6> CONF_DEC1<7>
                        + CONF_DEC1<8> CONF_DEC1<9> CONF_ROOUTFREQSEL<0> CONF_ROOUTFREQSEL<1>
                        + CONF_ROOUTFREQSEL<2> CONF_ROOUTFREQSEL<3> CONF_ROOUTSEL<0>
                        + CONF_ROOUTSEL<1> CONF_SELDC<0> CONF_SELDC<1> CONF_SELTDC<0> CONF_SELTDC<1>
                        + CONF_SENDFREE CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2>
                        + CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6>
                        + CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10>
                        + CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14>
                        + CONF_STATECNT<15> CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2>
                        + CONF_TDC00N<3> CONF_TDC00N<4> CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7>
                        + CONF_TDC00N<8> CONF_TDC00N<9> CONF_TDC00N<10> CONF_TDC00N<11>
                        + CONF_TDC00N<12> CONF_TDC00N<13> CONF_TDC00N<14> CONF_TDC00N<15>
                        + CONF_TDC00N<16> CONF_TDC00N<17> CONF_TDC00N<18> CONF_TDC00N<19>
                        + CONF_TDC00P<0> CONF_TDC00P<1> CONF_TDC00P<2> CONF_TDC00P<3> CONF_TDC00P<4>
                        + CONF_TDC00P<5> CONF_TDC00P<6> CONF_TDC00P<7> CONF_TDC00P<8> CONF_TDC00P<9>
                        + CONF_TDC00P<10> CONF_TDC00P<11> CONF_TDC00P<12> CONF_TDC00P<13>
                        + CONF_TDC00P<14> CONF_TDC00P<15> CONF_TDC00P<16> CONF_TDC00P<17>
                        + CONF_TDC00P<18> CONF_TDC00P<19> CONF_TDC01N<0> CONF_TDC01N<1>
                        + CONF_TDC01N<2> CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5> CONF_TDC01N<6>
                        + CONF_TDC01N<7> CONF_TDC01N<8> CONF_TDC01N<9> CONF_TDC01N<10>
                        + CONF_TDC01N<11> CONF_TDC01N<12> CONF_TDC01N<13> CONF_TDC01N<14>
                        + CONF_TDC01N<15> CONF_TDC01N<16> CONF_TDC01N<17> CONF_TDC01N<18>
                        + CONF_TDC01N<19> CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2>
                        + CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5> CONF_TDC01P<6> CONF_TDC01P<7>
                        + CONF_TDC01P<8> CONF_TDC01P<9> CONF_TDC01P<10> CONF_TDC01P<11>
                        + CONF_TDC01P<12> CONF_TDC01P<13> CONF_TDC01P<14> CONF_TDC01P<15>
                        + CONF_TDC01P<16> CONF_TDC01P<17> CONF_TDC01P<18> CONF_TDC01P<19> CONF_TDC4B
                        + CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2> CONF_TDC10N<3> CONF_TDC10N<4>
                        + CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10N<8> CONF_TDC10N<9>
                        + CONF_TDC10N<10> CONF_TDC10N<11> CONF_TDC10N<12> CONF_TDC10N<13>
                        + CONF_TDC10N<14> CONF_TDC10N<15> CONF_TDC10N<16> CONF_TDC10N<17>
                        + CONF_TDC10N<18> CONF_TDC10N<19> CONF_TDC10P<0> CONF_TDC10P<1>
                        + CONF_TDC10P<2> CONF_TDC10P<3> CONF_TDC10P<4> CONF_TDC10P<5> CONF_TDC10P<6>
                        + CONF_TDC10P<7> CONF_TDC10P<8> CONF_TDC10P<9> CONF_TDC10P<10>
                        + CONF_TDC10P<11> CONF_TDC10P<12> CONF_TDC10P<13> CONF_TDC10P<14>
                        + CONF_TDC10P<15> CONF_TDC10P<16> CONF_TDC10P<17> CONF_TDC10P<18>
                        + CONF_TDC10P<19> CONF_TDC11N<0> CONF_TDC11N<1> CONF_TDC11N<2>
                        + CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5> CONF_TDC11N<6> CONF_TDC11N<7>
                        + CONF_TDC11N<8> CONF_TDC11N<9> CONF_TDC11N<10> CONF_TDC11N<11>
                        + CONF_TDC11N<12> CONF_TDC11N<13> CONF_TDC11N<14> CONF_TDC11N<15>
                        + CONF_TDC11N<16> CONF_TDC11N<17> CONF_TDC11N<18> CONF_TDC11N<19>
                        + CONF_TDC11P<0> CONF_TDC11P<1> CONF_TDC11P<2> CONF_TDC11P<3> CONF_TDC11P<4>
                        + CONF_TDC11P<5> CONF_TDC11P<6> CONF_TDC11P<7> CONF_TDC11P<8> CONF_TDC11P<9>
                        + CONF_TDC11P<10> CONF_TDC11P<11> CONF_TDC11P<12> CONF_TDC11P<13>
                        + CONF_TDC11P<14> CONF_TDC11P<15> CONF_TDC11P<16> CONF_TDC11P<17>
                        + CONF_TDC11P<18> CONF_TDC11P<19> CONF_TDCCAL<0> CONF_TDCCAL<1>
                        + CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4> CONF_TDCCAL<5> CONF_TDCCAL<6>
                        + CONF_TDCCAL<7> CONF_TDCCAL<8> CONF_TDCCAL<9> CONF_TDCCNT<0> CONF_TDCCNT<1>
                        + CONF_TDCCNT<2> CONF_TDCCNT<3> CONF_TDCCNT<4> CONF_TDCCNT<5> CONF_TDCCNT<6>
                        + CONF_TDCCNT<7> CONF_TDCCNT<8> CONF_TDCCNT<9> CONF_TDCCNT<10>
                        + CONF_TDCCNT<11> CONF_TDCCNT<12> CONF_TDCCNT<13> CONF_TDCCNT<14>
                        + CONF_TDCCNT<15> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2>
                        + CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7>
                        + CONF_TDCWAIT<0> CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3>
                        + CONF_TDCWAIT<4> CONF_TDCWAIT<5> CONF_TDCWAIT<6> CONF_TDCWAIT<7> DATA_OUT
                        + DATA_OUT_I<3> DATA_READY DATA_READY_I<3> ENABLE_E2L ENABLE_E2L_I<3>
                        + EXT_CLK RO_ENABLE RO_ENABLE_I<3> RO_OUT RST SCAN_OUT<0> SCAN_OUT<1>
                        + SCAN_OUT<2> SCAN_OUT<3> SCAN_OUT<4> SCAN_OUT<5> SCAN_OUT<6> SCAN_OUT<7>
                        + SCAN_OUT<8> SCAN_OUT<9> SCAN_OUT<10> SCAN_OUT<11> SCAN_OUT<12>
                        + SCAN_OUT<13> SCAN_OUT<14> SCAN_OUT<15> SCAN_OUT<16> SCAN_OUT<17>
                        + SCAN_OUT<18> SCAN_OUT<19> SCAN_OUT<20> SCAN_OUT<21> SCAN_OUT<22> SER_CLK
                        + TRNG_RST TRNG_RST'_I<3> TRNG_RST_I<3> VDD_CORE VDD_DC VDD_TDC VSS
    Xi0 ALARM0<0> ALARM0<1> ALARM1<0> ALARM1<1> ALARM_DC CLK CONF_DEC0<0> CONF_DEC0<1> CONF_DEC0<2>
        + CONF_DEC0<3> CONF_DEC0<4> CONF_DEC0<5> CONF_DEC0<6> CONF_DEC0<7> CONF_DEC0<8> CONF_DEC0<9>
        + CONF_DEC1<0> CONF_DEC1<1> CONF_DEC1<2> CONF_DEC1<3> CONF_DEC1<4> CONF_DEC1<5> CONF_DEC1<6>
        + CONF_DEC1<7> CONF_DEC1<8> CONF_DEC1<9> CONF_SELDC<0> CONF_SELDC<1> CONF_SELTDC<0>
        + CONF_SELTDC<1> CONF_TDC00N<0> CONF_TDC00N<1> CONF_TDC00N<2> CONF_TDC00N<3> CONF_TDC00N<4>
        + CONF_TDC00N<5> CONF_TDC00N<6> CONF_TDC00N<7> CONF_TDC00N<8> CONF_TDC00N<9> CONF_TDC00N<10>
        + CONF_TDC00N<11> CONF_TDC00N<12> CONF_TDC00N<13> CONF_TDC00N<14> CONF_TDC00N<15>
        + CONF_TDC00N<16> CONF_TDC00N<17> CONF_TDC00N<18> CONF_TDC00N<19> CONF_TDC00P<0>
        + CONF_TDC00P<1> CONF_TDC00P<2> CONF_TDC00P<3> CONF_TDC00P<4> CONF_TDC00P<5> CONF_TDC00P<6>
        + CONF_TDC00P<7> CONF_TDC00P<8> CONF_TDC00P<9> CONF_TDC00P<10> CONF_TDC00P<11>
        + CONF_TDC00P<12> CONF_TDC00P<13> CONF_TDC00P<14> CONF_TDC00P<15> CONF_TDC00P<16>
        + CONF_TDC00P<17> CONF_TDC00P<18> CONF_TDC00P<19> CONF_TDC01N<0> CONF_TDC01N<1>
        + CONF_TDC01N<2> CONF_TDC01N<3> CONF_TDC01N<4> CONF_TDC01N<5> CONF_TDC01N<6> CONF_TDC01N<7>
        + CONF_TDC01N<8> CONF_TDC01N<9> CONF_TDC01N<10> CONF_TDC01N<11> CONF_TDC01N<12>
        + CONF_TDC01N<13> CONF_TDC01N<14> CONF_TDC01N<15> CONF_TDC01N<16> CONF_TDC01N<17>
        + CONF_TDC01N<18> CONF_TDC01N<19> CONF_TDC01P<0> CONF_TDC01P<1> CONF_TDC01P<2>
        + CONF_TDC01P<3> CONF_TDC01P<4> CONF_TDC01P<5> CONF_TDC01P<6> CONF_TDC01P<7> CONF_TDC01P<8>
        + CONF_TDC01P<9> CONF_TDC01P<10> CONF_TDC01P<11> CONF_TDC01P<12> CONF_TDC01P<13>
        + CONF_TDC01P<14> CONF_TDC01P<15> CONF_TDC01P<16> CONF_TDC01P<17> CONF_TDC01P<18>
        + CONF_TDC01P<19> CONF_TDC4B CONF_TDC10N<0> CONF_TDC10N<1> CONF_TDC10N<2> CONF_TDC10N<3>
        + CONF_TDC10N<4> CONF_TDC10N<5> CONF_TDC10N<6> CONF_TDC10N<7> CONF_TDC10N<8> CONF_TDC10N<9>
        + CONF_TDC10N<10> CONF_TDC10N<11> CONF_TDC10N<12> CONF_TDC10N<13> CONF_TDC10N<14>
        + CONF_TDC10N<15> CONF_TDC10N<16> CONF_TDC10N<17> CONF_TDC10N<18> CONF_TDC10N<19>
        + CONF_TDC10P<0> CONF_TDC10P<1> CONF_TDC10P<2> CONF_TDC10P<3> CONF_TDC10P<4> CONF_TDC10P<5>
        + CONF_TDC10P<6> CONF_TDC10P<7> CONF_TDC10P<8> CONF_TDC10P<9> CONF_TDC10P<10>
        + CONF_TDC10P<11> CONF_TDC10P<12> CONF_TDC10P<13> CONF_TDC10P<14> CONF_TDC10P<15>
        + CONF_TDC10P<16> CONF_TDC10P<17> CONF_TDC10P<18> CONF_TDC10P<19> CONF_TDC11N<0>
        + CONF_TDC11N<1> CONF_TDC11N<2> CONF_TDC11N<3> CONF_TDC11N<4> CONF_TDC11N<5> CONF_TDC11N<6>
        + CONF_TDC11N<7> CONF_TDC11N<8> CONF_TDC11N<9> CONF_TDC11N<10> CONF_TDC11N<11>
        + CONF_TDC11N<12> CONF_TDC11N<13> CONF_TDC11N<14> CONF_TDC11N<15> CONF_TDC11N<16>
        + CONF_TDC11N<17> CONF_TDC11N<18> CONF_TDC11N<19> CONF_TDC11P<0> CONF_TDC11P<1>
        + CONF_TDC11P<2> CONF_TDC11P<3> CONF_TDC11P<4> CONF_TDC11P<5> CONF_TDC11P<6> CONF_TDC11P<7>
        + CONF_TDC11P<8> CONF_TDC11P<9> CONF_TDC11P<10> CONF_TDC11P<11> CONF_TDC11P<12>
        + CONF_TDC11P<13> CONF_TDC11P<14> CONF_TDC11P<15> CONF_TDC11P<16> CONF_TDC11P<17>
        + CONF_TDC11P<18> CONF_TDC11P<19> CONF_TDCMAX<0> CONF_TDCMAX<1> CONF_TDCMAX<2>
        + CONF_TDCMAX<3> CONF_TDCMAX<4> CONF_TDCMAX<5> CONF_TDCMAX<6> CONF_TDCMAX<7> CONF_TDCWAIT<0>
        + CONF_TDCWAIT<1> CONF_TDCWAIT<2> CONF_TDCWAIT<3> CONF_TDCWAIT<4> CONF_TDCWAIT<5>
        + CONF_TDCWAIT<6> CONF_TDCWAIT<7> DCEDGE0<1> DCEDGE0<2> DCEDGE0<3> DCEDGE1<1> DCEDGE1<2>
        + DCEDGE1<3> DCEDGE2<1> DCEDGE2<2> DCEDGE2<3> ENABLE_E2L RO_ENABLE FF0<0> FF0<1> FF0<2>
        + FF0<3> FF0<4> FF0<5> FF0<6> FF0<7> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF1<5> FF1<6> FF1<7>
        + INT0 INT1 RO_OUT_I<0> RO_OUT_I<1> RO_OUT_I<2> RAND0 RAND1 READY0 READY1 TRNG_RST TRNG_RST'
        + CONF_DCEDGESEL<0> CONF_DCEDGESEL<1> SENDFREE'<8> SENDFREE'<9> SENDFREE'<16> SENDFREE'<0>
        + SENDFREE'<1> SENDFREE'<12> SENDFREE'<2> SENDFREE'<3> SENDFREE'<13> SENDFREE'<10>
        + SENDFREE'<11> SENDFREE'<17> SENDFREE'<4> SENDFREE'<5> SENDFREE'<14> SENDFREE'<6>
        + SENDFREE'<7> SENDFREE'<15> VDD_CORE VDD_DC VDD_TDC VSS trng_toplevel
    Xi1 ENABLE_E2L_I<0> CAL_OUT0 CAL_OUT1 CAL_OUT2 RO_OUT_I<3> RO_ENABLE_I<0> CLK CONF_STATECNT<0>
        + CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5>
        + CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10>
        + CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15>
        + CONF_TDCCAL<0> CONF_TDCCAL<1> CONF_TDCCAL<2> CONF_TDCCAL<3> CONF_TDCCAL<4> CONF_TDCCAL<5>
        + CONF_TDCCAL<6> CONF_TDCCAL<7> CONF_TDCCAL<8> CONF_TDCCAL<9> DATA_OUT_I<0> DATA_READY_I<0>
        + TRNG_RST_I<0> TRNG_RST'_I<0> RST_I RST'_I SER_CLK SCAN_OUT<3> SCAN_OUT<0> SCAN_OUT<1>
        + SCAN_OUT<2> SCAN_OUT<5> ALARM0<0> ALARM0<1> FF0<0> FF0<1> FF0<2> FF0<3> FF0<4> FF0<5>
        + FF0<6> FF0<7> INT0 READY0 ALARM1<0> ALARM1<1> FF1<0> FF1<1> FF1<2> FF1<3> FF1<4> FF1<5>
        + FF1<6> FF1<7> INT1 READY1 SCAN_OUT<4> VDD_CORE VSS conf_toplevel
    Xi2 ALARM_DC CLK CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2> CONF_STATECNT<3>
        + CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7> CONF_STATECNT<8>
        + CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12> CONF_STATECNT<13>
        + CONF_STATECNT<14> CONF_STATECNT<15> DATA_OUT_I<1> DATA_READY_I<1> TRNG_RST_I<1>
        + TRNG_RST'_I<1> RO_OUT_I<1> ENABLE_E2L_I<1> RO_ENABLE_I<1> RAND0 RAND1 RST_I RST'_I
        + CONF_SENDFREE SER_CLK SCAN_OUT<9> SCAN_OUT<6> SCAN_OUT<7> SCAN_OUT<8> SCAN_OUT<11>
        + ALARM0<0> ALARM0<1> READY0 ALARM1<0> ALARM1<1> READY1 SCAN_OUT<10> VDD_CORE VSS
        + bit_toplevel
    Xi3 CLK SCAN_OUT<17> SCAN_OUT<21> CONF_STATECNT<0> CONF_STATECNT<1> CONF_STATECNT<2>
        + CONF_STATECNT<3> CONF_STATECNT<4> CONF_STATECNT<5> CONF_STATECNT<6> CONF_STATECNT<7>
        + CONF_STATECNT<8> CONF_STATECNT<9> CONF_STATECNT<10> CONF_STATECNT<11> CONF_STATECNT<12>
        + CONF_STATECNT<13> CONF_STATECNT<14> CONF_STATECNT<15> CONF_TDCCNT<0> CONF_TDCCNT<1>
        + CONF_TDCCNT<2> CONF_TDCCNT<3> CONF_TDCCNT<4> CONF_TDCCNT<5> CONF_TDCCNT<6> CONF_TDCCNT<7>
        + CONF_TDCCNT<8> CONF_TDCCNT<9> CONF_TDCCNT<10> CONF_TDCCNT<11> CONF_TDCCNT<12>
        + CONF_TDCCNT<13> CONF_TDCCNT<14> CONF_TDCCNT<15> DATA_OUT_I<2> DATA_READY_I<2>
        + TRNG_RST_I<2> TRNG_RST'_I<2> SCAN_OUT<18> ENABLE_E2L_I<2> RO_ENABLE_I<2> RST_I RST'_I
        + SER_CLK SCAN_OUT<22> SCAN_OUT<12> SCAN_OUT<13> SCAN_OUT<14> SCAN_OUT<15> SCAN_OUT<16>
        + SCAN_OUT<20> READY0 READY1 SCAN_OUT<19> VDD_CORE VSS async_toplevel
    Xi26 RO_OUT_I<0> RO_OUT_I<1> RO_OUT_I<2> RO_OUT_I<3> RO_OUT_SEL CONF_ROOUTSEL<0>
         + CONF_ROOUTSEL<1> VDD_CORE VSS mux4
    Xi15 RO_ENABLE_I<0> RO_ENABLE_I<1> RO_ENABLE_I<2> RO_ENABLE_I<3> net028 CONF_CTRLSEL<0>
         + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi13 ENABLE_E2L_I<0> ENABLE_E2L_I<1> ENABLE_E2L_I<2> ENABLE_E2L_I<3> net024 CONF_CTRLSEL<0>
         + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi11 DATA_READY_I<0> DATA_READY_I<1> DATA_READY_I<2> DATA_READY_I<3> net0162 CONF_CTRLSEL<0>
         + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi9 DATA_OUT_I<0> DATA_OUT_I<1> DATA_OUT_I<2> DATA_OUT_I<3> net012 CONF_CTRLSEL<0>
        + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi5 TRNG_RST'_I<0> TRNG_RST'_I<1> TRNG_RST'_I<2> TRNG_RST'_I<3> net0157 CONF_CTRLSEL<0>
        + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi4 TRNG_RST_I<0> TRNG_RST_I<1> TRNG_RST_I<2> TRNG_RST_I<3> net0149 CONF_CTRLSEL<0>
        + CONF_CTRLSEL<1> VDD_CORE VSS mux4
    Xi36 net073 CLK VDD_CORE VSS buffer_large
    Xi33 RST RST_I VDD_CORE VSS buffer_large
    Xi32 RST' RST'_I VDD_CORE VSS buffer_large
    Xi30 net0142 RO_OUT VDD_CORE VSS buffer_large
    Xi16 net028 RO_ENABLE VDD_CORE VSS buffer_large
    Xi14 net024 ENABLE_E2L VDD_CORE VSS buffer_large
    Xi12 net0162 DATA_READY VDD_CORE VSS buffer_large
    Xi10 net012 DATA_OUT VDD_CORE VSS buffer_large
    Xi7 net0157 TRNG_RST' VDD_CORE VSS buffer_large
    Xi6 net0149 TRNG_RST VDD_CORE VSS buffer_large
    Xi25 CAL_OUT2 DCEDGE2<1> VDD_CORE VSS buffer
    Xi24 CAL_OUT1 DCEDGE2<3> VDD_CORE VSS buffer
    Xi23 CAL_OUT0 DCEDGE2<2> VDD_CORE VSS buffer
    Xi22 CAL_OUT2 DCEDGE1<2> VDD_CORE VSS buffer
    Xi21 CAL_OUT1 DCEDGE1<1> VDD_CORE VSS buffer
    Xi20 CAL_OUT0 DCEDGE1<3> VDD_CORE VSS buffer
    Xi19 CAL_OUT2 DCEDGE0<3> VDD_CORE VSS buffer
    Xi18 CAL_OUT1 DCEDGE0<2> VDD_CORE VSS buffer
    Xi17 CAL_OUT0 DCEDGE0<1> VDD_CORE VSS buffer
    Xi28 RO_OUT_SEL ROOUTFreq<0> ROOUTFreq<1> ROOUTFreq<2> ROOUTFreq<3> ROOUTFreq<4> ROOUTFreq<5>
         + ROOUTFreq<6> ROOUTFreq<7> ROOUTFreq<8> ROOUTFreq<9> ROOUTFreq<10> ROOUTFreq<11>
         + ROOUTFreq<12> ROOUTFreq<13> ROOUTFreq<14> ROOUTFreq<15> net0138 RST_I RST'_I VDD_CORE VSS
         + freq_scaler16
    Xi29 ROOUTFreq<0> ROOUTFreq<1> ROOUTFreq<2> ROOUTFreq<3> ROOUTFreq<4> ROOUTFreq<5> ROOUTFreq<6>
         + ROOUTFreq<7> ROOUTFreq<8> ROOUTFreq<9> ROOUTFreq<10> ROOUTFreq<11> ROOUTFreq<12>
         + ROOUTFreq<13> ROOUTFreq<14> ROOUTFreq<15> net0142 CONF_ROOUTFREQSEL<0>
         + CONF_ROOUTFREQSEL<1> CONF_ROOUTFREQSEL<2> CONF_ROOUTFREQSEL<3> VDD_CORE VSS mux16
    Xi31 RST RST' VDD_CORE VSS inv
    Xi34 GEN_CLK CONF_CLK<0> CONF_CLK<1> CONF_CLK<2> CONF_CLK<3> CONF_CLK<4> CONF_CLK<5> CONF_CLK<6>
         + CONF_CLK<7> CONF_CLK<8> CONF_CLK<9> CONF_CLK<10> CONF_CLK<11> CONF_CLKENABLE RST_I RST'_I
         + VDD_CORE VSS clkmanager
    Xi35 GEN_CLK EXT_CLK net073 CONF_CLKSEL VDD_CORE VSS mux2
    Xi37 CONF_SENDFREE SENDFREE'<0> SENDFREE'<1> SENDFREE'<2> SENDFREE'<3> SENDFREE'<4> SENDFREE'<5>
         + SENDFREE'<6> SENDFREE'<7> SENDFREE'<8> SENDFREE'<9> SENDFREE'<10> SENDFREE'<11>
         + SENDFREE'<12> SENDFREE'<13> SENDFREE'<14> SENDFREE'<15> SENDFREE'<16> SENDFREE'<17>
         + VDD_CORE VSS oneto18
.ENDS

.SUBCKT oneto7 IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> VDD VSS
    Xi6 IN OUT<6> VDD VSS inv
    Xi5 IN OUT<3> VDD VSS inv
    Xi4 IN OUT<5> VDD VSS inv
    Xi3 IN OUT<4> VDD VSS inv
    Xi2 IN OUT<2> VDD VSS inv
    Xi1 IN OUT<1> VDD VSS inv
    Xi0 IN OUT<0> VDD VSS inv
.ENDS

.SUBCKT conf_2 CLK IN OUT<0> OUT<1> RST RST' VDD VSS
    Xi1 CLK OUT<0> OUT<1> net14 RST RST' VDD VSS dff_st_ar_buf
    Xi0 CLK IN OUT<0> net13 RST RST' VDD VSS dff_st_ar_buf
.ENDS

.SUBCKT conf_4 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS
    Xi1 CLK OUT<1> OUT<2> OUT<3> RST RST' VDD VSS conf_2
    Xi0 CLK IN OUT<0> OUT<1> RST RST' VDD VSS conf_2
.ENDS

.SUBCKT conf_8 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS
    Xi1 CLK OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS conf_4
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS conf_4
.ENDS

.SUBCKT conf_16 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
                + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
    Xi1 CLK OUT<7> OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
        + conf_8
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS conf_8
.ENDS

.SUBCKT conf_32 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
                + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20>
                + OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30>
                + OUT<31> RST RST' VDD VSS
    Xi1 CLK OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25>
        + OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST' VDD VSS conf_16
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10> OUT<11>
        + OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS conf_16
.ENDS

.SUBCKT conf_64 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
                + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20>
                + OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30>
                + OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40>
                + OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50>
                + OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60>
                + OUT<61> OUT<62> OUT<63> RST RST' VDD VSS
    Xi1 CLK OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41>
        + OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52>
        + OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63>
        + RST RST' VDD VSS conf_32
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10> OUT<11>
        + OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22>
        + OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST' VDD VSS
        + conf_32
.ENDS

.SUBCKT conf_128 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                 + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                 + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                 + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                 + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                 + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                 + OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69>
                 + OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79>
                 + OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88> OUT<89>
                 + OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
                 + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107> OUT<108>
                 + OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115> OUT<116> OUT<117>
                 + OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125> OUT<126>
                 + OUT<127> RST RST' VDD VSS
    Xi1 CLK OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69> OUT<70> OUT<71> OUT<72> OUT<73>
        + OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79> OUT<80> OUT<81> OUT<82> OUT<83> OUT<84>
        + OUT<85> OUT<86> OUT<87> OUT<88> OUT<89> OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95>
        + OUT<96> OUT<97> OUT<98> OUT<99> OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105>
        + OUT<106> OUT<107> OUT<108> OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115>
        + OUT<116> OUT<117> OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125>
        + OUT<126> OUT<127> RST RST' VDD VSS conf_64
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10> OUT<11>
        + OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22>
        + OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32> OUT<33>
        + OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43> OUT<44>
        + OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55>
        + OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63> RST RST' VDD VSS conf_64
.ENDS

.SUBCKT conf_256 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                 + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                 + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                 + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                 + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                 + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                 + OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69>
                 + OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79>
                 + OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88> OUT<89>
                 + OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
                 + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107> OUT<108>
                 + OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115> OUT<116> OUT<117>
                 + OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125> OUT<126>
                 + OUT<127> OUT<128> OUT<129> OUT<130> OUT<131> OUT<132> OUT<133> OUT<134> OUT<135>
                 + OUT<136> OUT<137> OUT<138> OUT<139> OUT<140> OUT<141> OUT<142> OUT<143> OUT<144>
                 + OUT<145> OUT<146> OUT<147> OUT<148> OUT<149> OUT<150> OUT<151> OUT<152> OUT<153>
                 + OUT<154> OUT<155> OUT<156> OUT<157> OUT<158> OUT<159> OUT<160> OUT<161> OUT<162>
                 + OUT<163> OUT<164> OUT<165> OUT<166> OUT<167> OUT<168> OUT<169> OUT<170> OUT<171>
                 + OUT<172> OUT<173> OUT<174> OUT<175> OUT<176> OUT<177> OUT<178> OUT<179> OUT<180>
                 + OUT<181> OUT<182> OUT<183> OUT<184> OUT<185> OUT<186> OUT<187> OUT<188> OUT<189>
                 + OUT<190> OUT<191> OUT<192> OUT<193> OUT<194> OUT<195> OUT<196> OUT<197> OUT<198>
                 + OUT<199> OUT<200> OUT<201> OUT<202> OUT<203> OUT<204> OUT<205> OUT<206> OUT<207>
                 + OUT<208> OUT<209> OUT<210> OUT<211> OUT<212> OUT<213> OUT<214> OUT<215> OUT<216>
                 + OUT<217> OUT<218> OUT<219> OUT<220> OUT<221> OUT<222> OUT<223> OUT<224> OUT<225>
                 + OUT<226> OUT<227> OUT<228> OUT<229> OUT<230> OUT<231> OUT<232> OUT<233> OUT<234>
                 + OUT<235> OUT<236> OUT<237> OUT<238> OUT<239> OUT<240> OUT<241> OUT<242> OUT<243>
                 + OUT<244> OUT<245> OUT<246> OUT<247> OUT<248> OUT<249> OUT<250> OUT<251> OUT<252>
                 + OUT<253> OUT<254> OUT<255> RST RST' VDD VSS
    Xi1 CLK OUT<127> OUT<128> OUT<129> OUT<130> OUT<131> OUT<132> OUT<133> OUT<134> OUT<135>
        + OUT<136> OUT<137> OUT<138> OUT<139> OUT<140> OUT<141> OUT<142> OUT<143> OUT<144> OUT<145>
        + OUT<146> OUT<147> OUT<148> OUT<149> OUT<150> OUT<151> OUT<152> OUT<153> OUT<154> OUT<155>
        + OUT<156> OUT<157> OUT<158> OUT<159> OUT<160> OUT<161> OUT<162> OUT<163> OUT<164> OUT<165>
        + OUT<166> OUT<167> OUT<168> OUT<169> OUT<170> OUT<171> OUT<172> OUT<173> OUT<174> OUT<175>
        + OUT<176> OUT<177> OUT<178> OUT<179> OUT<180> OUT<181> OUT<182> OUT<183> OUT<184> OUT<185>
        + OUT<186> OUT<187> OUT<188> OUT<189> OUT<190> OUT<191> OUT<192> OUT<193> OUT<194> OUT<195>
        + OUT<196> OUT<197> OUT<198> OUT<199> OUT<200> OUT<201> OUT<202> OUT<203> OUT<204> OUT<205>
        + OUT<206> OUT<207> OUT<208> OUT<209> OUT<210> OUT<211> OUT<212> OUT<213> OUT<214> OUT<215>
        + OUT<216> OUT<217> OUT<218> OUT<219> OUT<220> OUT<221> OUT<222> OUT<223> OUT<224> OUT<225>
        + OUT<226> OUT<227> OUT<228> OUT<229> OUT<230> OUT<231> OUT<232> OUT<233> OUT<234> OUT<235>
        + OUT<236> OUT<237> OUT<238> OUT<239> OUT<240> OUT<241> OUT<242> OUT<243> OUT<244> OUT<245>
        + OUT<246> OUT<247> OUT<248> OUT<249> OUT<250> OUT<251> OUT<252> OUT<253> OUT<254> OUT<255>
        + RST RST' VDD VSS conf_128
    Xi0 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10> OUT<11>
        + OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22>
        + OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32> OUT<33>
        + OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43> OUT<44>
        + OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55>
        + OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66>
        + OUT<67> OUT<68> OUT<69> OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77>
        + OUT<78> OUT<79> OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88>
        + OUT<89> OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
        + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107> OUT<108> OUT<109>
        + OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115> OUT<116> OUT<117> OUT<118> OUT<119>
        + OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125> OUT<126> OUT<127> RST RST' VDD VSS
        + conf_128
.ENDS

.SUBCKT conf_268 CLK IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                 + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                 + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                 + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                 + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                 + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                 + OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69>
                 + OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79>
                 + OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88> OUT<89>
                 + OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
                 + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107> OUT<108>
                 + OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115> OUT<116> OUT<117>
                 + OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125> OUT<126>
                 + OUT<127> OUT<128> OUT<129> OUT<130> OUT<131> OUT<132> OUT<133> OUT<134> OUT<135>
                 + OUT<136> OUT<137> OUT<138> OUT<139> OUT<140> OUT<141> OUT<142> OUT<143> OUT<144>
                 + OUT<145> OUT<146> OUT<147> OUT<148> OUT<149> OUT<150> OUT<151> OUT<152> OUT<153>
                 + OUT<154> OUT<155> OUT<156> OUT<157> OUT<158> OUT<159> OUT<160> OUT<161> OUT<162>
                 + OUT<163> OUT<164> OUT<165> OUT<166> OUT<167> OUT<168> OUT<169> OUT<170> OUT<171>
                 + OUT<172> OUT<173> OUT<174> OUT<175> OUT<176> OUT<177> OUT<178> OUT<179> OUT<180>
                 + OUT<181> OUT<182> OUT<183> OUT<184> OUT<185> OUT<186> OUT<187> OUT<188> OUT<189>
                 + OUT<190> OUT<191> OUT<192> OUT<193> OUT<194> OUT<195> OUT<196> OUT<197> OUT<198>
                 + OUT<199> OUT<200> OUT<201> OUT<202> OUT<203> OUT<204> OUT<205> OUT<206> OUT<207>
                 + OUT<208> OUT<209> OUT<210> OUT<211> OUT<212> OUT<213> OUT<214> OUT<215> OUT<216>
                 + OUT<217> OUT<218> OUT<219> OUT<220> OUT<221> OUT<222> OUT<223> OUT<224> OUT<225>
                 + OUT<226> OUT<227> OUT<228> OUT<229> OUT<230> OUT<231> OUT<232> OUT<233> OUT<234>
                 + OUT<235> OUT<236> OUT<237> OUT<238> OUT<239> OUT<240> OUT<241> OUT<242> OUT<243>
                 + OUT<244> OUT<245> OUT<246> OUT<247> OUT<248> OUT<249> OUT<250> OUT<251> OUT<252>
                 + OUT<253> OUT<254> OUT<255> OUT<256> OUT<257> OUT<258> OUT<259> OUT<260> OUT<261>
                 + OUT<262> OUT<263> OUT<264> OUT<265> OUT<266> OUT<267> RST VDD VSS
    Xi0 CLK_I IN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21>
        + OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32>
        + OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43>
        + OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> OUT<53> OUT<54>
        + OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65>
        + OUT<66> OUT<67> OUT<68> OUT<69> OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76>
        + OUT<77> OUT<78> OUT<79> OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87>
        + OUT<88> OUT<89> OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98>
        + OUT<99> OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107> OUT<108>
        + OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115> OUT<116> OUT<117> OUT<118>
        + OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125> OUT<126> OUT<127> OUT<128>
        + OUT<129> OUT<130> OUT<131> OUT<132> OUT<133> OUT<134> OUT<135> OUT<136> OUT<137> OUT<138>
        + OUT<139> OUT<140> OUT<141> OUT<142> OUT<143> OUT<144> OUT<145> OUT<146> OUT<147> OUT<148>
        + OUT<149> OUT<150> OUT<151> OUT<152> OUT<153> OUT<154> OUT<155> OUT<156> OUT<157> OUT<158>
        + OUT<159> OUT<160> OUT<161> OUT<162> OUT<163> OUT<164> OUT<165> OUT<166> OUT<167> OUT<168>
        + OUT<169> OUT<170> OUT<171> OUT<172> OUT<173> OUT<174> OUT<175> OUT<176> OUT<177> OUT<178>
        + OUT<179> OUT<180> OUT<181> OUT<182> OUT<183> OUT<184> OUT<185> OUT<186> OUT<187> OUT<188>
        + OUT<189> OUT<190> OUT<191> OUT<192> OUT<193> OUT<194> OUT<195> OUT<196> OUT<197> OUT<198>
        + OUT<199> OUT<200> OUT<201> OUT<202> OUT<203> OUT<204> OUT<205> OUT<206> OUT<207> OUT<208>
        + OUT<209> OUT<210> OUT<211> OUT<212> OUT<213> OUT<214> OUT<215> OUT<216> OUT<217> OUT<218>
        + OUT<219> OUT<220> OUT<221> OUT<222> OUT<223> OUT<224> OUT<225> OUT<226> OUT<227> OUT<228>
        + OUT<229> OUT<230> OUT<231> OUT<232> OUT<233> OUT<234> OUT<235> OUT<236> OUT<237> OUT<238>
        + OUT<239> OUT<240> OUT<241> OUT<242> OUT<243> OUT<244> OUT<245> OUT<246> OUT<247> OUT<248>
        + OUT<249> OUT<250> OUT<251> OUT<252> OUT<253> OUT<254> OUT<255> RST_I RST'_I VDD VSS
        + conf_256
    Xi1 CLK_I OUT<255> OUT<256> OUT<257> OUT<258> OUT<259> OUT<260> OUT<261> OUT<262> OUT<263> RST_I
        + RST'_I VDD VSS conf_8
    Xi3 RST RST' VDD VSS inv
    Xi5 RST RST_I VDD VSS buffer_large
    Xi4 RST' RST'_I VDD VSS buffer_large
    Xi6 CLK CLK_I VDD VSS buffer_large
    Xi2 CLK_I OUT<263> OUT<264> OUT<265> OUT<266> OUT<267> RST_I RST'_I VDD VSS conf_4
.ENDS

.SUBCKT ctrl_trng_conf_combo CONF<260> CONF<261> CONF<262> CONF<263> CONF<264> CONF<265> CONF<266>
                             + CONF<267> CONF_CLK CONF_IN CONF_RST CORE_RST DATA_OUT DATA_READY
                             + EXT_CLK RO_OUT SCAN<0> SCAN<1> SCAN<2> SCAN<3> SCAN<4> SCAN<5>
                             + SCAN<6> SCAN<7> SCAN<8> SCAN<9> SCAN<10> SCAN<11> SCAN<12> SCAN<13>
                             + SCAN<14> SCAN<15> SCAN<16> SCAN<17> SCAN<18> SCAN<19> SCAN<20>
                             + SCAN<21> SCAN<22> SCAN<23> SCAN<24> SCAN<25> SENDFREE'<6> SER_CLK
                             + VDD_CORE VDD_DC VDD_TDC VSS
    Xi1 CONF<253> CONF<254> CONF<255> CONF<256> CONF<257> CONF<258> CONF<259> CONF<260> CONF<261>
        + CONF<262> CONF<263> CONF<264> CONF<265> CONF<252> CONF<0> CONF<1> CONF<49> CONF<50>
        + CONF<67> CONF<68> CONF<69> CONF<70> CONF<71> CONF<72> CONF<73> CONF<74> CONF<75> CONF<76>
        + CONF<77> CONF<78> CONF<79> CONF<80> CONF<81> CONF<82> CONF<83> CONF<84> CONF<85> CONF<86>
        + CONF<2> CONF<3> CONF<4> CONF<5> CONF<266> CONF<267> CONF<247> CONF<248> CONF<249>
        + CONF<250> CONF<48> CONF<16> CONF<17> CONF<18> CONF<19> CONF<20> CONF<21> CONF<22> CONF<23>
        + CONF<24> CONF<25> CONF<26> CONF<27> CONF<28> CONF<29> CONF<30> CONF<31> CONF<107>
        + CONF<108> CONF<109> CONF<110> CONF<111> CONF<112> CONF<113> CONF<114> CONF<115> CONF<116>
        + CONF<117> CONF<118> CONF<119> CONF<120> CONF<121> CONF<122> CONF<123> CONF<124> CONF<125>
        + CONF<126> CONF<87> CONF<88> CONF<89> CONF<90> CONF<91> CONF<92> CONF<93> CONF<94> CONF<95>
        + CONF<96> CONF<97> CONF<98> CONF<99> CONF<100> CONF<101> CONF<102> CONF<103> CONF<104>
        + CONF<105> CONF<106> CONF<147> CONF<148> CONF<149> CONF<150> CONF<151> CONF<152> CONF<153>
        + CONF<154> CONF<155> CONF<156> CONF<157> CONF<158> CONF<159> CONF<160> CONF<161> CONF<162>
        + CONF<163> CONF<164> CONF<165> CONF<166> CONF<127> CONF<128> CONF<129> CONF<130> CONF<131>
        + CONF<132> CONF<133> CONF<134> CONF<135> CONF<136> CONF<137> CONF<138> CONF<139> CONF<140>
        + CONF<141> CONF<142> CONF<143> CONF<144> CONF<145> CONF<146> CONF<251> CONF<187> CONF<188>
        + CONF<189> CONF<190> CONF<191> CONF<192> CONF<193> CONF<194> CONF<195> CONF<196> CONF<197>
        + CONF<198> CONF<199> CONF<200> CONF<201> CONF<202> CONF<203> CONF<204> CONF<205> CONF<206>
        + CONF<167> CONF<168> CONF<169> CONF<170> CONF<171> CONF<172> CONF<173> CONF<174> CONF<175>
        + CONF<176> CONF<177> CONF<178> CONF<179> CONF<180> CONF<181> CONF<182> CONF<183> CONF<184>
        + CONF<185> CONF<186> CONF<227> CONF<228> CONF<229> CONF<230> CONF<231> CONF<232> CONF<233>
        + CONF<234> CONF<235> CONF<236> CONF<237> CONF<238> CONF<239> CONF<240> CONF<241> CONF<242>
        + CONF<243> CONF<244> CONF<245> CONF<246> CONF<207> CONF<208> CONF<209> CONF<210> CONF<211>
        + CONF<212> CONF<213> CONF<214> CONF<215> CONF<216> CONF<217> CONF<218> CONF<219> CONF<220>
        + CONF<221> CONF<222> CONF<223> CONF<224> CONF<225> CONF<226> CONF<6> CONF<7> CONF<8>
        + CONF<9> CONF<10> CONF<11> CONF<12> CONF<13> CONF<14> CONF<15> CONF<32> CONF<33> CONF<34>
        + CONF<35> CONF<36> CONF<37> CONF<38> CONF<39> CONF<40> CONF<41> CONF<42> CONF<43> CONF<44>
        + CONF<45> CONF<46> CONF<47> CONF<59> CONF<60> CONF<61> CONF<62> CONF<63> CONF<64> CONF<65>
        + CONF<66> CONF<51> CONF<52> CONF<53> CONF<54> CONF<55> CONF<56> CONF<57> CONF<58> DATA_OUT
        + SENDFREE'<2> DATA_READY SENDFREE'<3> SCAN<25> SENDFREE'<4> EXT_CLK SCAN<24> SENDFREE'<5>
        + RO_OUT CORE_RST SCAN<0> SCAN<1> SCAN<2> SCAN<3> SCAN<4> SCAN<5> SCAN<6> SCAN<7> SCAN<8>
        + SCAN<9> SCAN<10> SCAN<11> SCAN<12> SCAN<13> SCAN<14> SCAN<15> SCAN<16> SCAN<17> SCAN<18>
        + SCAN<19> SCAN<20> SCAN<21> SCAN<22> SER_CLK SCAN<23> SENDFREE'<1> SENDFREE'<0> VDD_CORE
        + VDD_DC VDD_TDC VSS ctrl_trng_combo
    Xi2 CONF<48> SENDFREE'<0> SENDFREE'<1> SENDFREE'<2> SENDFREE'<3> SENDFREE'<4> SENDFREE'<5>
        + SENDFREE'<6> VDD_CORE VSS oneto7
    Xi0 CONF_CLK CONF_IN CONF<0> CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> CONF<8>
        + CONF<9> CONF<10> CONF<11> CONF<12> CONF<13> CONF<14> CONF<15> CONF<16> CONF<17> CONF<18>
        + CONF<19> CONF<20> CONF<21> CONF<22> CONF<23> CONF<24> CONF<25> CONF<26> CONF<27> CONF<28>
        + CONF<29> CONF<30> CONF<31> CONF<32> CONF<33> CONF<34> CONF<35> CONF<36> CONF<37> CONF<38>
        + CONF<39> CONF<40> CONF<41> CONF<42> CONF<43> CONF<44> CONF<45> CONF<46> CONF<47> CONF<48>
        + CONF<49> CONF<50> CONF<51> CONF<52> CONF<53> CONF<54> CONF<55> CONF<56> CONF<57> CONF<58>
        + CONF<59> CONF<60> CONF<61> CONF<62> CONF<63> CONF<64> CONF<65> CONF<66> CONF<67> CONF<68>
        + CONF<69> CONF<70> CONF<71> CONF<72> CONF<73> CONF<74> CONF<75> CONF<76> CONF<77> CONF<78>
        + CONF<79> CONF<80> CONF<81> CONF<82> CONF<83> CONF<84> CONF<85> CONF<86> CONF<87> CONF<88>
        + CONF<89> CONF<90> CONF<91> CONF<92> CONF<93> CONF<94> CONF<95> CONF<96> CONF<97> CONF<98>
        + CONF<99> CONF<100> CONF<101> CONF<102> CONF<103> CONF<104> CONF<105> CONF<106> CONF<107>
        + CONF<108> CONF<109> CONF<110> CONF<111> CONF<112> CONF<113> CONF<114> CONF<115> CONF<116>
        + CONF<117> CONF<118> CONF<119> CONF<120> CONF<121> CONF<122> CONF<123> CONF<124> CONF<125>
        + CONF<126> CONF<127> CONF<128> CONF<129> CONF<130> CONF<131> CONF<132> CONF<133> CONF<134>
        + CONF<135> CONF<136> CONF<137> CONF<138> CONF<139> CONF<140> CONF<141> CONF<142> CONF<143>
        + CONF<144> CONF<145> CONF<146> CONF<147> CONF<148> CONF<149> CONF<150> CONF<151> CONF<152>
        + CONF<153> CONF<154> CONF<155> CONF<156> CONF<157> CONF<158> CONF<159> CONF<160> CONF<161>
        + CONF<162> CONF<163> CONF<164> CONF<165> CONF<166> CONF<167> CONF<168> CONF<169> CONF<170>
        + CONF<171> CONF<172> CONF<173> CONF<174> CONF<175> CONF<176> CONF<177> CONF<178> CONF<179>
        + CONF<180> CONF<181> CONF<182> CONF<183> CONF<184> CONF<185> CONF<186> CONF<187> CONF<188>
        + CONF<189> CONF<190> CONF<191> CONF<192> CONF<193> CONF<194> CONF<195> CONF<196> CONF<197>
        + CONF<198> CONF<199> CONF<200> CONF<201> CONF<202> CONF<203> CONF<204> CONF<205> CONF<206>
        + CONF<207> CONF<208> CONF<209> CONF<210> CONF<211> CONF<212> CONF<213> CONF<214> CONF<215>
        + CONF<216> CONF<217> CONF<218> CONF<219> CONF<220> CONF<221> CONF<222> CONF<223> CONF<224>
        + CONF<225> CONF<226> CONF<227> CONF<228> CONF<229> CONF<230> CONF<231> CONF<232> CONF<233>
        + CONF<234> CONF<235> CONF<236> CONF<237> CONF<238> CONF<239> CONF<240> CONF<241> CONF<242>
        + CONF<243> CONF<244> CONF<245> CONF<246> CONF<247> CONF<248> CONF<249> CONF<250> CONF<251>
        + CONF<252> CONF<253> CONF<254> CONF<255> CONF<256> CONF<257> CONF<258> CONF<259> CONF<260>
        + CONF<261> CONF<262> CONF<263> CONF<264> CONF<265> CONF<266> CONF<267> CONF_RST VDD_CORE
        + VSS conf_268
.ENDS

.SUBCKT scan_1 CLK IN_PAR IN_SER OUT RST RST' SER VDD VSS
    Xi0 IN_PAR IN_SER net19 SER VDD VSS mux2
    Xi1 CLK net19 OUT net21 RST RST' VDD VSS dff_st_ar
.ENDS

.SUBCKT scan_2 CLK IN_PAR<0> IN_PAR<1> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK IN_PAR<1> net13 OUT RST RST' SER VDD VSS scan_1
    Xi0 CLK IN_PAR<0> IN_SER net13 RST RST' SER VDD VSS scan_1
.ENDS

.SUBCKT scan_4 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK IN_PAR<2> IN_PAR<3> net13 OUT RST RST' SER VDD VSS scan_2
    Xi0 CLK IN_PAR<0> IN_PAR<1> IN_SER net13 RST RST' SER VDD VSS scan_2
.ENDS

.SUBCKT scan_8 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
               + IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> net13 OUT RST RST' SER VDD VSS scan_4
    Xi0 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER net13 RST RST' SER VDD VSS scan_4
.ENDS

.SUBCKT scan_16 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
                + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14>
                + IN_PAR<15> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + net13 OUT RST RST' SER VDD VSS scan_8
    Xi0 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> IN_SER
        + net13 RST RST' SER VDD VSS scan_8
.ENDS

.SUBCKT scan_32 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
                + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14>
                + IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21>
                + IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28>
                + IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + net13 OUT RST RST' SER VDD VSS scan_16
    Xi0 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_SER net13 RST RST' SER VDD VSS scan_16
.ENDS

.SUBCKT scan_34 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
                + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14>
                + IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21>
                + IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28>
                + IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_PAR<32> IN_PAR<33> IN_SER OUT RST SER VDD VSS
    Xi2 RST RST' VDD VSS inv
    Xi0 CLK_I IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + IN_SER net13 RST_I RST'_I SER_I VDD VSS scan_32
    Xi1 CLK_I IN_PAR<32> IN_PAR<33> net13 OUT_I RST_I RST'_I SER_I VDD VSS scan_2
    Xi7 OUT_I OUT VDD VSS buffer_large
    Xi6 SER SER_I VDD VSS buffer_large
    Xi5 CLK CLK_I VDD VSS buffer_large
    Xi4 RST RST_I VDD VSS buffer_large
    Xi3 RST' RST'_I VDD VSS buffer_large
.ENDS

.SUBCKT ctrl_trng_conf_scan_combo CONF_CLK CONF_IN CONF_RST CORE_RST DATA_OUT DATA_READY EXT_CLK
                                  + RO_OUT SCAN_CLK SCAN_OUT SCAN_RST SCAN_SER SER_CLK VDD_CORE
                                  + VDD_DC VDD_TDC VSS
    Xi0 SCAN<26> SCAN<27> SCAN<28> SCAN<29> SCAN<30> SCAN<31> SCAN<32> SCAN<33> CONF_CLK CONF_IN
        + CONF_RST CORE_RST DATA_OUT DATA_READY EXT_CLK RO_OUT SCAN<0> SCAN<1> SCAN<2> SCAN<3>
        + SCAN<4> SCAN<5> SCAN<6> SCAN<7> SCAN<8> SCAN<9> SCAN<10> SCAN<11> SCAN<12> SCAN<13>
        + SCAN<14> SCAN<15> SCAN<16> SCAN<17> SCAN<18> SCAN<19> SCAN<20> SCAN<21> SCAN<22> SCAN<23>
        + SCAN<24> SCAN<25> net21 SER_CLK VDD_CORE VDD_DC VDD_TDC VSS ctrl_trng_conf_combo
    Xi1 SCAN_CLK SCAN<0> SCAN<1> SCAN<2> SCAN<3> SCAN<4> SCAN<5> SCAN<6> SCAN<7> SCAN<8> SCAN<9>
        + SCAN<10> SCAN<11> SCAN<12> SCAN<13> SCAN<14> SCAN<15> SCAN<16> SCAN<17> SCAN<18> SCAN<19>
        + SCAN<20> SCAN<21> SCAN<22> SCAN<23> SCAN<24> SCAN<25> SCAN<26> SCAN<27> SCAN<28> SCAN<29>
        + SCAN<30> SCAN<31> SCAN<32> SCAN<33> net21 SCAN_OUT SCAN_RST SCAN_SER VDD_CORE VSS scan_34
.ENDS

.SUBCKT inv_jit IN OUT VDD VSS
    Mm0 OUT IN VDD VDD p_mos l=60n w=480.0n m=1
    Mm1 OUT IN VSS VSS n_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dc_jit_2 CLK IN LAST OUT<0> OUT<1> RST RST' VDD VSS
    Xi3 CLK LAST OUT<1> net24 RST RST' VDD VSS dff_st_ar
    Xi2 CLK INT net25 OUT<0> RST RST' VDD VSS dff_st_ar
    Xi1 INT LAST VDD VSS inv_jit
    Xi0 IN INT VDD VSS inv_jit
.ENDS

.SUBCKT dc_jit_4 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<2> OUT<3> RST RST' VDD VSS dc_jit_2
    Xi0 CLK IN INT OUT<0> OUT<1> RST RST' VDD VSS dc_jit_2
.ENDS

.SUBCKT dc_jit_8 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD
                 + VSS
    Xi1 CLK INT LAST OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS dc_jit_4
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS dc_jit_4
.ENDS

.SUBCKT dc_jit_16 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
        + dc_jit_8
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS dc_jit_8
.ENDS

.SUBCKT dc_jit_32 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                  + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                  + OUT<30> OUT<31> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25>
        + OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST' VDD VSS dc_jit_16
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS dc_jit_16
.ENDS

.SUBCKT dc_jit_64 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                  + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                  + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                  + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                  + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                  + OUT<60> OUT<61> OUT<62> OUT<63> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41>
        + OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52>
        + OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63>
        + RST RST' VDD VSS dc_jit_32
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21>
        + OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST'
        + VDD VSS dc_jit_32
.ENDS

.SUBCKT dc_jit_128 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                   + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                   + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                   + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                   + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                   + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                   + OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69>
                   + OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79>
                   + OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88> OUT<89>
                   + OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
                   + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107>
                   + OUT<108> OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115>
                   + OUT<116> OUT<117> OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123>
                   + OUT<124> OUT<125> OUT<126> OUT<127> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69> OUT<70> OUT<71> OUT<72> OUT<73>
        + OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79> OUT<80> OUT<81> OUT<82> OUT<83> OUT<84>
        + OUT<85> OUT<86> OUT<87> OUT<88> OUT<89> OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95>
        + OUT<96> OUT<97> OUT<98> OUT<99> OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105>
        + OUT<106> OUT<107> OUT<108> OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115>
        + OUT<116> OUT<117> OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125>
        + OUT<126> OUT<127> RST RST' VDD VSS dc_jit_64
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21>
        + OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32>
        + OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43>
        + OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> OUT<53> OUT<54>
        + OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63> RST RST' VDD VSS
        + dc_jit_64
.ENDS

.SUBCKT scan_jit_2 CLK IN_PAR<0> IN_PAR<1> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK net12 OUT net14 RST RST' VDD VSS dff_st_ar
    Xi0 CLK net07 net11 net15 RST RST' VDD VSS dff_st_ar
    Xi4 IN_PAR<0> IN_SER net07 SER VDD VSS mux2
    Xi2 IN_PAR<1> net11 net12 SER VDD VSS mux2
.ENDS

.SUBCKT scan_jit_4 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_SER net8 RST RST' SER VDD VSS scan_jit_2
    Xi6 CLK IN_PAR<2> IN_PAR<3> net8 OUT RST RST' SER VDD VSS scan_jit_2
.ENDS

.SUBCKT scan_jit_8 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                   + IN_PAR<7> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER net8 RST RST' SER VDD VSS scan_jit_4
    Xi6 CLK IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> net8 OUT RST RST' SER VDD VSS scan_jit_4
.ENDS

.SUBCKT scan_jit_16 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> IN_SER
        + net8 RST RST' SER VDD VSS scan_jit_8
    Xi6 CLK IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + net8 OUT RST RST' SER VDD VSS scan_jit_8
.ENDS

.SUBCKT scan_jit_32 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                    + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                    + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_16
    Xi6 CLK IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + net8 OUT RST RST' SER VDD VSS scan_jit_16
.ENDS

.SUBCKT scan_jit_64 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                    + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                    + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_PAR<32> IN_PAR<33> IN_PAR<34>
                    + IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39> IN_PAR<40> IN_PAR<41>
                    + IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47> IN_PAR<48>
                    + IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
                    + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62>
                    + IN_PAR<63> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_32
    Xi6 CLK IN_PAR<32> IN_PAR<33> IN_PAR<34> IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39>
        + IN_PAR<40> IN_PAR<41> IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47>
        + IN_PAR<48> IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
        + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62> IN_PAR<63>
        + net8 OUT RST RST' SER VDD VSS scan_jit_32
.ENDS

.SUBCKT scan_jit_128 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                     + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                     + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                     + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                     + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_PAR<32> IN_PAR<33> IN_PAR<34>
                     + IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39> IN_PAR<40> IN_PAR<41>
                     + IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47> IN_PAR<48>
                     + IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
                     + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62>
                     + IN_PAR<63> IN_PAR<64> IN_PAR<65> IN_PAR<66> IN_PAR<67> IN_PAR<68> IN_PAR<69>
                     + IN_PAR<70> IN_PAR<71> IN_PAR<72> IN_PAR<73> IN_PAR<74> IN_PAR<75> IN_PAR<76>
                     + IN_PAR<77> IN_PAR<78> IN_PAR<79> IN_PAR<80> IN_PAR<81> IN_PAR<82> IN_PAR<83>
                     + IN_PAR<84> IN_PAR<85> IN_PAR<86> IN_PAR<87> IN_PAR<88> IN_PAR<89> IN_PAR<90>
                     + IN_PAR<91> IN_PAR<92> IN_PAR<93> IN_PAR<94> IN_PAR<95> IN_PAR<96> IN_PAR<97>
                     + IN_PAR<98> IN_PAR<99> IN_PAR<100> IN_PAR<101> IN_PAR<102> IN_PAR<103>
                     + IN_PAR<104> IN_PAR<105> IN_PAR<106> IN_PAR<107> IN_PAR<108> IN_PAR<109>
                     + IN_PAR<110> IN_PAR<111> IN_PAR<112> IN_PAR<113> IN_PAR<114> IN_PAR<115>
                     + IN_PAR<116> IN_PAR<117> IN_PAR<118> IN_PAR<119> IN_PAR<120> IN_PAR<121>
                     + IN_PAR<122> IN_PAR<123> IN_PAR<124> IN_PAR<125> IN_PAR<126> IN_PAR<127>
                     + IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + IN_PAR<32> IN_PAR<33> IN_PAR<34> IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39>
        + IN_PAR<40> IN_PAR<41> IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47>
        + IN_PAR<48> IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
        + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62> IN_PAR<63>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_64
    Xi6 CLK IN_PAR<64> IN_PAR<65> IN_PAR<66> IN_PAR<67> IN_PAR<68> IN_PAR<69> IN_PAR<70> IN_PAR<71>
        + IN_PAR<72> IN_PAR<73> IN_PAR<74> IN_PAR<75> IN_PAR<76> IN_PAR<77> IN_PAR<78> IN_PAR<79>
        + IN_PAR<80> IN_PAR<81> IN_PAR<82> IN_PAR<83> IN_PAR<84> IN_PAR<85> IN_PAR<86> IN_PAR<87>
        + IN_PAR<88> IN_PAR<89> IN_PAR<90> IN_PAR<91> IN_PAR<92> IN_PAR<93> IN_PAR<94> IN_PAR<95>
        + IN_PAR<96> IN_PAR<97> IN_PAR<98> IN_PAR<99> IN_PAR<100> IN_PAR<101> IN_PAR<102>
        + IN_PAR<103> IN_PAR<104> IN_PAR<105> IN_PAR<106> IN_PAR<107> IN_PAR<108> IN_PAR<109>
        + IN_PAR<110> IN_PAR<111> IN_PAR<112> IN_PAR<113> IN_PAR<114> IN_PAR<115> IN_PAR<116>
        + IN_PAR<117> IN_PAR<118> IN_PAR<119> IN_PAR<120> IN_PAR<121> IN_PAR<122> IN_PAR<123>
        + IN_PAR<124> IN_PAR<125> IN_PAR<126> IN_PAR<127> net8 OUT RST RST' SER VDD VSS scan_jit_64
.ENDS

.SUBCKT dc_scan_jit_128 DC_CLK DC_IN DC_LAST DC_RST DC_RST' SCAN_CLK SCAN_IN_SER SCAN_OUT SCAN_RST
                        + SCAN_RST' SCAN_SER VDD VSS
    Xi0 DC_CLK DC_IN DC_LAST DC_OUT<0> DC_OUT<1> DC_OUT<2> DC_OUT<3> DC_OUT<4> DC_OUT<5> DC_OUT<6>
        + DC_OUT<7> DC_OUT<8> DC_OUT<9> DC_OUT<10> DC_OUT<11> DC_OUT<12> DC_OUT<13> DC_OUT<14>
        + DC_OUT<15> DC_OUT<16> DC_OUT<17> DC_OUT<18> DC_OUT<19> DC_OUT<20> DC_OUT<21> DC_OUT<22>
        + DC_OUT<23> DC_OUT<24> DC_OUT<25> DC_OUT<26> DC_OUT<27> DC_OUT<28> DC_OUT<29> DC_OUT<30>
        + DC_OUT<31> DC_OUT<32> DC_OUT<33> DC_OUT<34> DC_OUT<35> DC_OUT<36> DC_OUT<37> DC_OUT<38>
        + DC_OUT<39> DC_OUT<40> DC_OUT<41> DC_OUT<42> DC_OUT<43> DC_OUT<44> DC_OUT<45> DC_OUT<46>
        + DC_OUT<47> DC_OUT<48> DC_OUT<49> DC_OUT<50> DC_OUT<51> DC_OUT<52> DC_OUT<53> DC_OUT<54>
        + DC_OUT<55> DC_OUT<56> DC_OUT<57> DC_OUT<58> DC_OUT<59> DC_OUT<60> DC_OUT<61> DC_OUT<62>
        + DC_OUT<63> DC_OUT<64> DC_OUT<65> DC_OUT<66> DC_OUT<67> DC_OUT<68> DC_OUT<69> DC_OUT<70>
        + DC_OUT<71> DC_OUT<72> DC_OUT<73> DC_OUT<74> DC_OUT<75> DC_OUT<76> DC_OUT<77> DC_OUT<78>
        + DC_OUT<79> DC_OUT<80> DC_OUT<81> DC_OUT<82> DC_OUT<83> DC_OUT<84> DC_OUT<85> DC_OUT<86>
        + DC_OUT<87> DC_OUT<88> DC_OUT<89> DC_OUT<90> DC_OUT<91> DC_OUT<92> DC_OUT<93> DC_OUT<94>
        + DC_OUT<95> DC_OUT<96> DC_OUT<97> DC_OUT<98> DC_OUT<99> DC_OUT<100> DC_OUT<101> DC_OUT<102>
        + DC_OUT<103> DC_OUT<104> DC_OUT<105> DC_OUT<106> DC_OUT<107> DC_OUT<108> DC_OUT<109>
        + DC_OUT<110> DC_OUT<111> DC_OUT<112> DC_OUT<113> DC_OUT<114> DC_OUT<115> DC_OUT<116>
        + DC_OUT<117> DC_OUT<118> DC_OUT<119> DC_OUT<120> DC_OUT<121> DC_OUT<122> DC_OUT<123>
        + DC_OUT<124> DC_OUT<125> DC_OUT<126> DC_OUT<127> DC_RST DC_RST' VDD VSS dc_jit_128
    Xi1 SCAN_CLK DC_OUT<0> DC_OUT<1> DC_OUT<2> DC_OUT<3> DC_OUT<4> DC_OUT<5> DC_OUT<6> DC_OUT<7>
        + DC_OUT<8> DC_OUT<9> DC_OUT<10> DC_OUT<11> DC_OUT<12> DC_OUT<13> DC_OUT<14> DC_OUT<15>
        + DC_OUT<16> DC_OUT<17> DC_OUT<18> DC_OUT<19> DC_OUT<20> DC_OUT<21> DC_OUT<22> DC_OUT<23>
        + DC_OUT<24> DC_OUT<25> DC_OUT<26> DC_OUT<27> DC_OUT<28> DC_OUT<29> DC_OUT<30> DC_OUT<31>
        + DC_OUT<32> DC_OUT<33> DC_OUT<34> DC_OUT<35> DC_OUT<36> DC_OUT<37> DC_OUT<38> DC_OUT<39>
        + DC_OUT<40> DC_OUT<41> DC_OUT<42> DC_OUT<43> DC_OUT<44> DC_OUT<45> DC_OUT<46> DC_OUT<47>
        + DC_OUT<48> DC_OUT<49> DC_OUT<50> DC_OUT<51> DC_OUT<52> DC_OUT<53> DC_OUT<54> DC_OUT<55>
        + DC_OUT<56> DC_OUT<57> DC_OUT<58> DC_OUT<59> DC_OUT<60> DC_OUT<61> DC_OUT<62> DC_OUT<63>
        + DC_OUT<64> DC_OUT<65> DC_OUT<66> DC_OUT<67> DC_OUT<68> DC_OUT<69> DC_OUT<70> DC_OUT<71>
        + DC_OUT<72> DC_OUT<73> DC_OUT<74> DC_OUT<75> DC_OUT<76> DC_OUT<77> DC_OUT<78> DC_OUT<79>
        + DC_OUT<80> DC_OUT<81> DC_OUT<82> DC_OUT<83> DC_OUT<84> DC_OUT<85> DC_OUT<86> DC_OUT<87>
        + DC_OUT<88> DC_OUT<89> DC_OUT<90> DC_OUT<91> DC_OUT<92> DC_OUT<93> DC_OUT<94> DC_OUT<95>
        + DC_OUT<96> DC_OUT<97> DC_OUT<98> DC_OUT<99> DC_OUT<100> DC_OUT<101> DC_OUT<102>
        + DC_OUT<103> DC_OUT<104> DC_OUT<105> DC_OUT<106> DC_OUT<107> DC_OUT<108> DC_OUT<109>
        + DC_OUT<110> DC_OUT<111> DC_OUT<112> DC_OUT<113> DC_OUT<114> DC_OUT<115> DC_OUT<116>
        + DC_OUT<117> DC_OUT<118> DC_OUT<119> DC_OUT<120> DC_OUT<121> DC_OUT<122> DC_OUT<123>
        + DC_OUT<124> DC_OUT<125> DC_OUT<126> DC_OUT<127> SCAN_IN_SER SCAN_OUT SCAN_RST SCAN_RST'
        + SCAN_SER VDD VSS scan_jit_128
.ENDS

.SUBCKT jit_top_half CONF<15> CONF_CLK CONF_IN CONF_RST CONF_RST' CORE_RST CORE_RST' DC_CLK
                     + RO_ENABLE RO_OUT SCAN_CLK SCAN_IN_SER SCAN_OUT SCAN_RST SCAN_RST' SCAN_SER
                     + VDD_CORE VDD_JIT VSS
    Xi0 RO CONF<0> CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> CONF<8> CONF<9> CONF<10>
        + CONF<11> RO_ENABLE CORE_RST CORE_RST' VDD_JIT VSS clkmanager
    Xi1 DC_CLK RO LAST CORE_RST CORE_RST' SCAN_CLK SCAN_IN_SER SCAN_INT SCAN_RST SCAN_RST' SCAN_SER
        + VDD_CORE VSS dc_scan_jit_128
    Xi2 CNT_CLK CNT<0> CNT<1> CNT<2> CNT<3> CNT<4> CNT<5> CNT<6> CNT<7> CNT<8> CNT<9> CNT<10>
        + CNT<11> CNT<12> CNT<13> CNT<14> CNT<15> CNT<16> CNT<17> CNT<18> CNT<19> CNT<20> CNT<21>
        + CNT<22> CNT<23> CNT<24> CNT<25> CNT<26> CNT<27> CNT<28> CNT<29> CNT<30> CNT<31> net22
        + CORE_RST CORE_RST' VDD_CORE VSS asynccounter_32
    Xi3 CNT<8> CNT<9> CNT<10> CNT<11> CNT<12> CNT<13> CNT<14> CNT<15> CNT<16> CNT<17> CNT<18>
        + CNT<19> CNT<20> CNT<21> CNT<22> CNT<23> RO_OUT_I CONF<12> CONF<13> CONF<14> CONF<15>
        + VDD_CORE VSS mux16
    Xi4 CONF_CLK CONF_IN CONF<0> CONF<1> CONF<2> CONF<3> CONF<4> CONF<5> CONF<6> CONF<7> CONF<8>
        + CONF<9> CONF<10> CONF<11> CONF<12> CONF<13> CONF<14> CONF<15> CONF_RST CONF_RST' VDD_CORE
        + VSS conf_16
    Xi5 SCAN_CLK CNT<0> CNT<1> CNT<2> CNT<3> CNT<4> CNT<5> CNT<6> CNT<7> CNT<8> CNT<9> CNT<10>
        + CNT<11> CNT<12> CNT<13> CNT<14> CNT<15> CNT<16> CNT<17> CNT<18> CNT<19> CNT<20> CNT<21>
        + CNT<22> CNT<23> CNT<24> CNT<25> CNT<26> CNT<27> CNT<28> CNT<29> CNT<30> CNT<31> SCAN_INT
        + SCAN_OUT_I SCAN_RST SCAN_RST' SCAN_SER VDD_CORE VSS scan_32
    Xi7 SCAN_OUT_I SCAN_OUT VDD_CORE VSS buffer_large
    Xi6 RO_OUT_I RO_OUT VDD_CORE VSS buffer_large
    Xi8 LAST DC_CLK CNT_CLK VDD_CORE VSS nor2
.ENDS

.SUBCKT jit_top_full CONF_CLK CONF_IN CONF_RST CORE_RST DC_CLK RO_ENABLE RO_OUT0 RO_OUT1 SCAN_CLK
                     + SCAN_OUT SCAN_RST SCAN_SER VDD_CORE VDD_JIT0 VDD_JIT1 VSS
    Xi1 net034 CONF_CLK_I CONF_INT CONF_RST_I CONF_RST'_I CORE_RST_I CORE_RST'_I DC_CLK_I RO_ENABLE
        + RO_OUT1 SCAN_CLK_I SCAN_OUT_INT SCAN_OUT SCAN_RST_I SCAN_RST'_I SCAN_SER_I VDD_CORE
        + VDD_JIT1 VSS jit_top_half
    Xi0 CONF_INT CONF_CLK_I CONF_IN CONF_RST_I CONF_RST'_I CORE_RST_I CORE_RST'_I DC_CLK_I RO_ENABLE
        + RO_OUT0 SCAN_CLK_I SCAN_OUT SCAN_OUT_INT SCAN_RST_I SCAN_RST'_I SCAN_SER_I VDD_CORE
        + VDD_JIT0 VSS jit_top_half
    Xi4 SCAN_RST SCAN_RST' VDD_CORE VSS inv
    Xi3 CONF_RST CONF_RST' VDD_CORE VSS inv
    Xi2 CORE_RST CORE_RST' VDD_CORE VSS inv
    Xi14 DC_CLK DC_CLK_I VDD_CORE VSS buffer_large
    Xi13 CONF_CLK CONF_CLK_I VDD_CORE VSS buffer_large
    Xi12 SCAN_CLK SCAN_CLK_I VDD_CORE VSS buffer_large
    Xi11 SCAN_SER SCAN_SER_I VDD_CORE VSS buffer_large
    Xi10 SCAN_RST SCAN_RST_I VDD_CORE VSS buffer_large
    Xi9 SCAN_RST' SCAN_RST'_I VDD_CORE VSS buffer_large
    Xi8 CONF_RST' CONF_RST'_I VDD_CORE VSS buffer_large
    Xi7 CONF_RST CONF_RST_I VDD_CORE VSS buffer_large
    Xi6 CORE_RST CORE_RST_I VDD_CORE VSS buffer_large
    Xi5 CORE_RST' CORE_RST'_I VDD_CORE VSS buffer_large
.ENDS

.SUBCKT top_core JIT_CONF_CLK JIT_CONF_IN JIT_CONF_RST JIT_CORE_RST JIT_DC_CLK JIT_RO_ENABLE
                 + JIT_RO_OUT0 JIT_RO_OUT1 JIT_SCAN_CLK JIT_SCAN_OUT JIT_SCAN_RST JIT_SCAN_SER
                 + JIT_VDD_CORE JIT_VDD_JIT0 JIT_VDD_JIT1 TRNG_CONF_CLK TRNG_CONF_IN TRNG_CONF_RST
                 + TRNG_CORE_RST TRNG_DATA_OUT TRNG_DATA_READY TRNG_EXT_CLK TRNG_RO_OUT
                 + TRNG_SCAN_CLK TRNG_SCAN_OUT TRNG_SCAN_RST TRNG_SCAN_SER TRNG_SER_CLK
                 + TRNG_VDD_CORE TRNG_VDD_DC TRNG_VDD_TDC VSS
    Xi0 TRNG_CONF_CLK TRNG_CONF_IN TRNG_CONF_RST TRNG_CORE_RST TRNG_DATA_OUT TRNG_DATA_READY
        + TRNG_EXT_CLK TRNG_RO_OUT TRNG_SCAN_CLK TRNG_SCAN_OUT TRNG_SCAN_RST TRNG_SCAN_SER
        + TRNG_SER_CLK TRNG_VDD_CORE TRNG_VDD_DC TRNG_VDD_TDC VSS ctrl_trng_conf_scan_combo
    Xi1 JIT_CONF_CLK JIT_CONF_IN JIT_CONF_RST JIT_CORE_RST JIT_DC_CLK JIT_RO_ENABLE JIT_RO_OUT0
        + JIT_RO_OUT1 JIT_SCAN_CLK JIT_SCAN_OUT JIT_SCAN_RST JIT_SCAN_SER JIT_VDD_CORE JIT_VDD_JIT0
        + JIT_VDD_JIT1 VSS jit_top_full
.ENDS

.SUBCKT decouplecap VDD VSS
    Mc0 VDD VSS VSS VSS cap nv=32 nh=32 w=100n s=100n stm=1 spm=4 m=300
.ENDS

.SUBCKT top_level JIT_CONF_CLK_PAD JIT_CONF_IN_PAD JIT_CONF_RST_PAD JIT_CORE_RST_PAD JIT_DC_CLK_PAD
                  + JIT_RO_ENABLE_PAD JIT_RO_OUT0_PAD JIT_RO_OUT1_PAD JIT_SCAN_CLK_PAD
                  + JIT_SCAN_OUT_PAD JIT_SCAN_RST_PAD JIT_SCAN_SER_PAD JIT_VDD_CORE_PAD
                  + JIT_VDD_JIT0_PAD JIT_VDD_JIT1_PAD TRNG_CONF_CLK_PAD TRNG_CONF_IN_PAD
                  + TRNG_CONF_RST_PAD TRNG_CORE_RST_PAD TRNG_DATA_OUT_PAD TRNG_DATA_READY_PAD
                  + TRNG_EXT_CLK_PAD TRNG_RO_OUT_PAD TRNG_SCAN_CLK_PAD TRNG_SCAN_OUT_PAD
                  + TRNG_SCAN_RST_PAD TRNG_SCAN_SER_PAD TRNG_SER_CLK_PAD TRNG_VDD_CORE_PAD
                  + TRNG_VDD_DC_PAD TRNG_VDD_TDC_PAD VDD_IO_PAD VSS_PAD
    Xi0 JIT_CONF_CLK JIT_CONF_CLK_PAD JIT_CONF_IN JIT_CONF_IN_PAD JIT_CONF_RST JIT_CONF_RST_PAD
        + JIT_CORE_RST JIT_CORE_RST_PAD JIT_DC_CLK JIT_DC_CLK_PAD JIT_RO_ENABLE JIT_RO_ENABLE_PAD
        + JIT_RO_OUT0 JIT_RO_OUT0_PAD JIT_RO_OUT1 JIT_RO_OUT1_PAD JIT_SCAN_CLK JIT_SCAN_CLK_PAD
        + JIT_SCAN_OUT JIT_SCAN_OUT_PAD JIT_SCAN_RST JIT_SCAN_RST_PAD JIT_SCAN_SER JIT_SCAN_SER_PAD
        + JIT_VDD_CORE_PAD JIT_VDD_JIT0_PAD JIT_VDD_JIT1_PAD TRNG_CONF_CLK TRNG_CONF_CLK_PAD
        + TRNG_CONF_IN TRNG_CONF_IN_PAD TRNG_CONF_RST TRNG_CONF_RST_PAD TRNG_CORE_RST
        + TRNG_CORE_RST_PAD TRNG_DATA_OUT TRNG_DATA_OUT_PAD TRNG_DATA_READY TRNG_DATA_READY_PAD
        + TRNG_EXT_CLK TRNG_EXT_CLK_PAD TRNG_RO_OUT TRNG_RO_OUT_PAD TRNG_SCAN_CLK TRNG_SCAN_CLK_PAD
        + TRNG_SCAN_OUT TRNG_SCAN_OUT_PAD TRNG_SCAN_RST TRNG_SCAN_RST_PAD TRNG_SCAN_SER
        + TRNG_SCAN_SER_PAD TRNG_SER_CLK TRNG_SER_CLK_PAD TRNG_VDD_CORE_PAD TRNG_VDD_DC_PAD
        + TRNG_VDD_TDC_PAD VDD_IO_PAD VSS_PAD padframe_v1
    Xi1 JIT_CONF_CLK JIT_CONF_IN JIT_CONF_RST JIT_CORE_RST JIT_DC_CLK JIT_RO_ENABLE JIT_RO_OUT0
        + JIT_RO_OUT1 JIT_SCAN_CLK JIT_SCAN_OUT JIT_SCAN_RST JIT_SCAN_SER JIT_VDD_CORE_PAD
        + JIT_VDD_JIT0_PAD JIT_VDD_JIT1_PAD TRNG_CONF_CLK TRNG_CONF_IN TRNG_CONF_RST TRNG_CORE_RST
        + TRNG_DATA_OUT TRNG_DATA_READY TRNG_EXT_CLK TRNG_RO_OUT TRNG_SCAN_CLK TRNG_SCAN_OUT
        + TRNG_SCAN_RST TRNG_SCAN_SER TRNG_SER_CLK TRNG_VDD_CORE_PAD TRNG_VDD_DC_PAD
        + TRNG_VDD_TDC_PAD VSS_PAD top_core
    Xi7 JIT_VDD_CORE_PAD VSS_PAD decouplecap
    Xi6 JIT_VDD_JIT1_PAD VSS_PAD decouplecap
    Xi5 JIT_VDD_JIT0_PAD VSS_PAD decouplecap
    Xi4 TRNG_VDD_TDC_PAD VSS_PAD decouplecap
    Xi3 TRNG_VDD_DC_PAD VSS_PAD decouplecap
    Xi2 TRNG_VDD_CORE_PAD VSS_PAD decouplecap
.ENDS
