* Top cell name: tdc_1b_diff_branch

.SUBCKT inv_wn in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=240.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm5 net17 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm4 net18 in1 net17 vss n_mos l=60n w=360.0n m=1
    Mm3 out in0 net18 vss n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=60n w=360.0n m=1
    Mm2 net5 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm1 net16 in1 net5 vss n_mos l=60n w=360.0n m=1
    Mm0 out in0 net16 vss n_mos l=60n w=360.0n m=1
    Mm7 net32 rst vdd vdd p_mos l=60n w=480.0n m=1
    Mm6 out in2 net32 vdd p_mos l=60n w=480.0n m=1
    Mm5 out in1 net32 vdd p_mos l=60n w=480.0n m=1
    Mm4 out in0 net32 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
.ENDS

.SUBCKT nor2 in0 in1 out vdd vss
    Mm1 out in1 vss vss n_mos l=60n w=120.0n m=1
    Mm0 out in0 vss vss n_mos l=60n w=120.0n m=1
    Mm3 net7 in1 vdd vdd p_mos l=60n w=480.0n m=1
    Mm2 out in0 net7 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=120.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT tdc_and_diff in0_n in0_p in1_n in1_p out_n out_p vdd vss
    Mm3 net18 in1_p vss vss n_mos l=60n w=240.0n m=1
    Mm2 out_n in0_p net18 vss n_mos l=60n w=240.0n m=1
    Mm1 out_p in0_n vss vss n_mos l=60n w=120.0n m=1
    Mm0 out_p in1_n vss vss n_mos l=60n w=120.0n m=1
    Mm5 out_n out_p vdd vdd p_mos l=60n w=120.0n m=1
    Mm4 out_p out_n vdd vdd p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_buf_diff_np_4lin conf_n<0> conf_n<1> conf_n<2> conf_n<3> conf_p<0> conf_p<1> conf_p<2>
                             + conf_p<3> in_n in_p out_n out_p vdd vss
    Mm51 conf_n'<3> conf_n<3> vss vss n_mos l=60n w=120.0n m=1
    Mm50 conf_n'<2> conf_n<2> vss vss n_mos l=60n w=120.0n m=1
    Mm49 conf_n'<1> conf_n<1> vss vss n_mos l=60n w=120.0n m=1
    Mm48 conf_n'<0> conf_n<0> vss vss n_mos l=60n w=120.0n m=1
    Mm43 conf_p'<3> conf_p<3> vss vss n_mos l=60n w=120.0n m=1
    Mm42 conf_p'<2> conf_p<2> vss vss n_mos l=60n w=120.0n m=1
    Mm41 conf_p'<1> conf_p<1> vss vss n_mos l=60n w=120.0n m=1
    Mm40 conf_p'<0> conf_p<0> vss vss n_mos l=60n w=120.0n m=1
    Mm35 out_p in_n vss vss n_mos l=60n w=120.0n m=1
    Mm33 out_n in_p vss vss n_mos l=60n w=120.0n m=1
    Mm15 net49 conf_n<3> vss vss n_mos l=60n w=120.0n m=1
    Mm14 net52 conf_n<2> vss vss n_mos l=60n w=120.0n m=1
    Mm13 net53 conf_n<1> vss vss n_mos l=60n w=120.0n m=1
    Mm12 net56 conf_n<0> vss vss n_mos l=60n w=120.0n m=1
    Mm11 out_p out_n net49 vss n_mos l=60n w=120.0n m=1
    Mm10 out_p out_n net52 vss n_mos l=60n w=120.0n m=1
    Mm9 out_p out_n net53 vss n_mos l=60n w=120.0n m=1
    Mm8 out_p out_n net56 vss n_mos l=60n w=120.0n m=1
    Mm7 net57 conf_p<3> vss vss n_mos l=60n w=120.0n m=1
    Mm6 net60 conf_p<2> vss vss n_mos l=60n w=120.0n m=1
    Mm5 net61 conf_p<1> vss vss n_mos l=60n w=120.0n m=1
    Mm4 net64 conf_p<0> vss vss n_mos l=60n w=120.0n m=1
    Mm3 out_n out_p net57 vss n_mos l=60n w=120.0n m=1
    Mm2 out_n out_p net60 vss n_mos l=60n w=120.0n m=1
    Mm1 out_n out_p net61 vss n_mos l=60n w=120.0n m=1
    Mm0 out_n out_p net64 vss n_mos l=60n w=120.0n m=1
    Mm47 conf_n'<3> conf_n<3> vdd vdd p_mos l=60n w=120.0n m=1
    Mm46 conf_n'<2> conf_n<2> vdd vdd p_mos l=60n w=120.0n m=1
    Mm45 conf_n'<1> conf_n<1> vdd vdd p_mos l=60n w=120.0n m=1
    Mm44 conf_n'<0> conf_n<0> vdd vdd p_mos l=60n w=120.0n m=1
    Mm39 conf_p'<3> conf_p<3> vdd vdd p_mos l=60n w=120.0n m=1
    Mm38 conf_p'<2> conf_p<2> vdd vdd p_mos l=60n w=120.0n m=1
    Mm37 conf_p'<1> conf_p<1> vdd vdd p_mos l=60n w=120.0n m=1
    Mm36 conf_p'<0> conf_p<0> vdd vdd p_mos l=60n w=120.0n m=1
    Mm34 out_p in_n vdd vdd p_mos l=60n w=120.0n m=1
    Mm32 out_n in_p vdd vdd p_mos l=60n w=120.0n m=1
    Mm31 out_p out_n net50 vdd p_mos l=60n w=120.0n m=1
    Mm30 out_p out_n net51 vdd p_mos l=60n w=120.0n m=1
    Mm29 out_p out_n net54 vdd p_mos l=60n w=120.0n m=1
    Mm28 out_p out_n net55 vdd p_mos l=60n w=120.0n m=1
    Mm27 net50 conf_p'<3> vdd vdd p_mos l=60n w=120.0n m=1
    Mm26 net51 conf_p'<2> vdd vdd p_mos l=60n w=120.0n m=1
    Mm25 net54 conf_p'<1> vdd vdd p_mos l=60n w=120.0n m=1
    Mm24 net55 conf_p'<0> vdd vdd p_mos l=60n w=120.0n m=1
    Mm23 out_n out_p net58 vdd p_mos l=60n w=120.0n m=1
    Mm22 out_n out_p net59 vdd p_mos l=60n w=120.0n m=1
    Mm21 out_n out_p net62 vdd p_mos l=60n w=120.0n m=1
    Mm20 out_n out_p net63 vdd p_mos l=60n w=120.0n m=1
    Mm19 net58 conf_n'<3> vdd vdd p_mos l=60n w=120.0n m=1
    Mm18 net59 conf_n'<2> vdd vdd p_mos l=60n w=120.0n m=1
    Mm17 net62 conf_n'<1> vdd vdd p_mos l=60n w=120.0n m=1
    Mm16 net63 conf_n'<0> vdd vdd p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_inv in out vdd vss
    Mm0 out in vdd vdd p_mos l=60n w=120.0n m=1
    Mm1 out in vss vss n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT tdc_inv_wide in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=480.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT tdc_stage_diff_np_4lin_buf conf_n<0> conf_n<1> conf_n<2> conf_n<3> conf_p<0> conf_p<1>
                                   + conf_p<2> conf_p<3> in0_n in0_p in1_n in1_p out_buf_n out_buf_p
                                   + out_n out_p vdd vss
    Xi0 in0_n in0_p in1_n in1_p int_n int_p vdd vss tdc_and_diff
    Xi1 conf_n<0> conf_n<1> conf_n<2> conf_n<3> conf_p<0> conf_p<1> conf_p<2> conf_p<3> int_n int_p
        + out_n_i out_p_i vdd vss tdc_buf_diff_np_4lin
    Xi3 out_n out_buf_p vdd vss tdc_inv
    Xi2 out_p out_buf_n vdd vss tdc_inv
    Xi4 out_n_i out_p vdd vss tdc_inv_wide
    Xi5 out_p_i out_n vdd vss tdc_inv_wide
.ENDS

.SUBCKT tdc_2stage_diff_np_4lin_buf buf0_n buf0_p buf1_n buf1_p conf0_n<0> conf0_n<1> conf0_n<2>
                                    + conf0_n<3> conf0_p<0> conf0_p<1> conf0_p<2> conf0_p<3>
                                    + conf1_n<0> conf1_n<1> conf1_n<2> conf1_n<3> conf1_p<0>
                                    + conf1_p<1> conf1_p<2> conf1_p<3> ff0 ff1 in0_n in0_p in1_n
                                    + in1_p nand0_in nand0_out nand1_in nand1_out out0_n out0_p
                                    + out1_n out1_p rst rst' vdd vss
    Xi19 out_buf1_n buf1_n vdd vss inv_wn
    Xi16 out_buf0_p buf0_p vdd vss inv_wn
    Xi17 out_buf0_n buf0_n vdd vss inv_wn
    Xi18 out_buf1_p buf1_p vdd vss inv_wn
    Xi13 nor0 nand0 ff0 q0' rst rst' vdd vss dff_st_ar
    Xi12 nor1 nand1 ff1 q1' rst rst' vdd vss dff_st_ar
    Xi10 q0' enable0 nand0_out vdd vss nand2
    Xi11 q1' enable1 nand1_out vdd vss nand2
    Xi6 q1' out_buf0_n nand1 vdd vss nand2
    Xi7 q0' out_buf1_p nand0 vdd vss nand2
    Xi9 out_buf0_p nand0_in nor0 vdd vss nor2
    Xi8 out_buf1_n nand1_in nor1 vdd vss nor2
    Xi15 nand0_in enable0 vdd vss inv
    Xi14 nand1_in enable1 vdd vss inv
    Xi1 conf1_n<0> conf1_n<1> conf1_n<2> conf1_n<3> conf1_p<0> conf1_p<1> conf1_p<2> conf1_p<3>
        + in1_n in1_p nand1_in enable1 out_buf1_n out_buf1_p out1_n out1_p vdd vss
        + tdc_stage_diff_np_4lin_buf
    Xi0 conf0_n<0> conf0_n<1> conf0_n<2> conf0_n<3> conf0_p<0> conf0_p<1> conf0_p<2> conf0_p<3>
        + in0_n in0_p nand0_in enable0 out_buf0_n out_buf0_p out0_n out0_p vdd vss
        + tdc_stage_diff_np_4lin_buf
.ENDS

.SUBCKT tdc_stage_diff_np_4lin_switched_buf conf_n<0> conf_n<1> conf_n<2> conf_n<3> conf_p<0>
                                            + conf_p<1> conf_p<2> conf_p<3> in0_n in0_p in1_n in1_p
                                            + out_buf_n out_buf_p out_n out_p vdd vss
    Xi0 in0_n in0_p in1_n in1_p int_n int_p vdd vss tdc_and_diff
    Xi1 conf_n<0> conf_n<1> conf_n<2> conf_n<3> conf_p<0> conf_p<1> conf_p<2> conf_p<3> int_p int_n
        + out_n_i out_p_i vdd vss tdc_buf_diff_np_4lin
    Xi3 out_n out_buf_p vdd vss tdc_inv
    Xi2 out_p out_buf_n vdd vss tdc_inv
    Xi4 out_n_i out_p vdd vss tdc_inv_wide
    Xi5 out_p_i out_n vdd vss tdc_inv_wide
.ENDS

.SUBCKT tdc_2stage_diff_np_4lin_switched_buf buf0_n buf0_p buf1_n buf1_p conf0_n<0> conf0_n<1>
                                             + conf0_n<2> conf0_n<3> conf0_p<0> conf0_p<1>
                                             + conf0_p<2> conf0_p<3> conf1_n<0> conf1_n<1>
                                             + conf1_n<2> conf1_n<3> conf1_p<0> conf1_p<1>
                                             + conf1_p<2> conf1_p<3> edge0_n edge0_p edge1_n edge1_p
                                             + ff0 ff1 in0_n in0_p in1_n in1_p nand0_in nand0_out
                                             + nand1_in nand1_out out0_n out0_p out1_n out1_p rst
                                             + rst' vdd vss
    Xi15 nand1_in rst' net059 vdd vss nand2
    Xi14 nand0_in rst' net036 vdd vss nand2
    Xi11 q1' net059 nand1_out vdd vss nand2
    Xi10 q0' net036 nand0_out vdd vss nand2
    Xi4 q0' out_buf1_p nand0 vdd vss nand2
    Xi5 q1' out_buf0_n nand1 vdd vss nand2
    Xi6 out_buf0_p nand0_in nor0 vdd vss nor2
    Xi7 out_buf1_n nand1_in nor1 vdd vss nor2
    Xi8 nor0 nand0 ff0 q0' rst rst' vdd vss dff_st_ar
    Xi9 nor1 nand1 ff1 q1' rst rst' vdd vss dff_st_ar
    Xi19 out_buf1_n buf1_n vdd vss inv_wn
    Xi18 out_buf1_p buf1_p vdd vss inv_wn
    Xi17 out_buf0_n buf0_n vdd vss inv_wn
    Xi16 out_buf0_p buf0_p vdd vss inv_wn
    Xi1 conf1_n<0> conf1_n<1> conf1_n<2> conf1_n<3> conf1_p<0> conf1_p<1> conf1_p<2> conf1_p<3>
        + in1_n in1_p edge1_n edge1_p out_buf1_n out_buf1_p out1_n out1_p vdd vss
        + tdc_stage_diff_np_4lin_switched_buf
    Xi0 conf0_n<0> conf0_n<1> conf0_n<2> conf0_n<3> conf0_p<0> conf0_p<1> conf0_p<2> conf0_p<3>
        + in0_n in0_p edge0_n edge0_p out_buf0_n out_buf0_p out0_n out0_p vdd vss
        + tdc_stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT tdc_2e_1b_diff_np_4lin_buf buf0_n<0> buf0_n<1> buf0_p<0> buf0_p<1> buf1_n<0> buf1_n<1>
                                   + buf1_p<0> buf1_p<1> conf0_n<0> conf0_n<1> conf0_n<2> conf0_n<3>
                                   + conf0_n<4> conf0_n<5> conf0_n<6> conf0_n<7> conf0_p<0>
                                   + conf0_p<1> conf0_p<2> conf0_p<3> conf0_p<4> conf0_p<5>
                                   + conf0_p<6> conf0_p<7> conf1_n<0> conf1_n<1> conf1_n<2>
                                   + conf1_n<3> conf1_n<4> conf1_n<5> conf1_n<6> conf1_n<7>
                                   + conf1_p<0> conf1_p<1> conf1_p<2> conf1_p<3> conf1_p<4>
                                   + conf1_p<5> conf1_p<6> conf1_p<7> edge0_n edge0_p edge1_n
                                   + edge1_p ff0<0> ff0<1> ff1<0> ff1<1> rst rst' vdd vss
    Xi13 buf0_n<1> buf0_p<1> buf1_n<1> buf1_p<1> conf0_n<4> conf0_n<5> conf0_n<6> conf0_n<7>
         + conf0_p<4> conf0_p<5> conf0_p<6> conf0_p<7> conf1_n<4> conf1_n<5> conf1_n<6> conf1_n<7>
         + conf1_p<4> conf1_p<5> conf1_p<6> conf1_p<7> ff0<1> ff1<1> int0_n<0> int0_p<0> int1_n<0>
         + int1_p<0> nand0<0> nand0<1> nand1<0> nand1<1> int0_n<1> int0_p<1> int1_n<1> int1_p<1> rst
         + rst' vdd vss tdc_2stage_diff_np_4lin_buf
    Xi12 buf0_n<0> buf0_p<0> buf1_n<0> buf1_p<0> conf0_n<0> conf0_n<1> conf0_n<2> conf0_n<3>
         + conf0_p<0> conf0_p<1> conf0_p<2> conf0_p<3> conf1_n<0> conf1_n<1> conf1_n<2> conf1_n<3>
         + conf1_p<0> conf1_p<1> conf1_p<2> conf1_p<3> edge0_n edge0_p edge1_n edge1_p ff0<0> ff1<0>
         + int1_n<1> int1_p<1> int0_n<1> int0_p<1> nand1<1> nand0<0> nand0<1> nand1<0> int0_n<0>
         + int0_p<0> int1_n<0> int1_p<0> rst rst' vdd vss tdc_2stage_diff_np_4lin_switched_buf
.ENDS

.SUBCKT dec_stage conf_rand ff_in ff_prev out vdd vss
    Xi0 ff_in net3 vdd vss inv
    Xi1 ff_prev net3 net4 vdd vss nor2
    Xi2 net4 conf_rand out vdd vss nand2
.ENDS

.SUBCKT dec_4_conf_0 conf_dec<0> conf_dec<1> conf_dec<2> conf_dec<3> ff_in<0> ff_in<1> ff_in<2>
                     + ff_in<3> rand_out vdd vss
    Xi27 conf_dec<3> ff_in<3> ff_in<2> stage<3> vdd vss dec_stage
    Xi21 conf_dec<2> ff_in<2> ff_in<1> stage<2> vdd vss dec_stage
    Xi19 conf_dec<1> ff_in<1> ff_in<0> stage<1> vdd vss dec_stage
    Xi18 conf_dec<0> ff_in<0> ff_in<3> stage<0> vdd vss dec_stage
    Xi26 net026 net023 rand_out vdd vss nor2
    Xi25 stage<2> stage<3> net023 vdd vss nand2
    Xi24 stage<0> stage<1> net026 vdd vss nand2
.ENDS

.SUBCKT tff_st_ar clk q q' rst rst' vdd vss
    Xi0 clk q' q q' rst rst' vdd vss dff_st_ar
.ENDS

.SUBCKT async_counter_8 clk out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> q' rst rst' vdd
                        + vss
    Xi7 net4 out<4> net5 rst rst' vdd vss tff_st_ar
    Xi6 net6 out<6> net7 rst rst' vdd vss tff_st_ar
    Xi5 net7 out<7> q' rst rst' vdd vss tff_st_ar
    Xi4 net5 out<5> net6 rst rst' vdd vss tff_st_ar
    Xi3 net2 out<2> net3 rst rst' vdd vss tff_st_ar
    Xi2 net3 out<3> net4 rst rst' vdd vss tff_st_ar
    Xi1 net1 out<1> net2 rst rst' vdd vss tff_st_ar
    Xi0 clk out<0> net1 rst rst' vdd vss tff_st_ar
.ENDS

.SUBCKT nand4 in0 in1 in2 in3 out vdd vss
    Mm3 out in3 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm7 net21 in3 vss vss n_mos l=60n w=480.0n m=1
    Mm6 net22 in2 net21 vss n_mos l=60n w=480.0n m=1
    Mm5 net23 in1 net22 vss n_mos l=60n w=480.0n m=1
    Mm4 out in0 net23 vss n_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar_dh clk q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
    Xi6 n1 n3 vdd vss inv_wn
.ENDS

.SUBCKT max_ready conf_maxcycles<0> conf_maxcycles<1> conf_maxcycles<2> conf_maxcycles<3>
                  + conf_maxcycles<4> conf_maxcycles<5> conf_maxcycles<6> conf_maxcycles<7> int
                  + max_ready rst rst' vdd vss
    Xi0 int cnt<0> cnt<1> cnt<2> cnt<3> cnt<4> cnt<5> cnt<6> cnt<7> net020 rst rst' vdd vss
        + async_counter_8
    Xi8 cnt<7> conf_maxcycles<7> cnt_high<7> vdd vss nand2
    Xi7 cnt<6> conf_maxcycles<6> cnt_high<6> vdd vss nand2
    Xi6 cnt<5> conf_maxcycles<5> cnt_high<5> vdd vss nand2
    Xi5 cnt<4> conf_maxcycles<4> cnt_high<4> vdd vss nand2
    Xi4 cnt<3> conf_maxcycles<3> cnt_high<3> vdd vss nand2
    Xi3 cnt<2> conf_maxcycles<2> cnt_high<2> vdd vss nand2
    Xi2 cnt<1> conf_maxcycles<1> cnt_high<1> vdd vss nand2
    Xi1 cnt<0> conf_maxcycles<0> cnt_high<0> vdd vss nand2
    Xi10 cnt_high<4> cnt_high<5> cnt_high<6> cnt_high<7> net09 vdd vss nand4
    Xi9 cnt_high<0> cnt_high<1> cnt_high<2> cnt_high<3> net010 vdd vss nand4
    Xi11 net010 net09 net021 vdd vss nor2
    Xi12 net021 ready vdd vss inv
    Xi13 ready max_ready net018 rst rst' vdd vss dff_st_ar_dh
.ENDS

.SUBCKT nor4 in0 in1 in2 in3 out vdd vss
    Mm3 out in0 net7 vdd p_mos l=60n w=480.0n m=1
    Mm2 net7 in1 net6 vdd p_mos l=60n w=480.0n m=1
    Mm1 net6 in2 net5 vdd p_mos l=60n w=480.0n m=1
    Mm0 net5 in3 vdd vdd p_mos l=60n w=480.0n m=1
    Mm7 out in3 vss vss n_mos l=60n w=120.0n m=1
    Mm6 out in2 vss vss n_mos l=60n w=120.0n m=1
    Mm5 out in0 vss vss n_mos l=60n w=120.0n m=1
    Mm4 out in1 vss vss n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT buffer in out vdd vss
    Mm1 out int vss vss n_mos l=60n w=480.0n m=4
    Mm0 int in vss vss n_mos l=60n w=480.0n m=1
    Mm3 out int vdd vdd p_mos l=60n w=480.0n m=4
    Mm2 int in vdd vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT wait_ready clk conf_waitcycles<0> conf_waitcycles<1> conf_waitcycles<2> conf_waitcycles<3>
                   + conf_waitcycles<4> conf_waitcycles<5> conf_waitcycles<6> conf_waitcycles<7>
                   + enable_e2l int rst rst' vdd vss wait_ready
    Xi4 clk_int wait_cnt<0> wait_cnt<1> wait_cnt<2> wait_cnt<3> wait_cnt<4> wait_cnt<5> wait_cnt<6>
        + wait_cnt<7> net044 cnt_rst cnt_rst' vdd vss async_counter_8
    Xi26 clk net049 net052 vdd vss nand2
    Xi19 wait_cnt<7> conf_waitcycles<7> waithigh<7> vdd vss nand2
    Xi18 wait_cnt<6> conf_waitcycles<6> waithigh<6> vdd vss nand2
    Xi17 wait_cnt<5> conf_waitcycles<5> waithigh<5> vdd vss nand2
    Xi10 wait_cnt<4> conf_waitcycles<4> waithigh<4> vdd vss nand2
    Xi3 wait_cnt<3> conf_waitcycles<3> waithigh<3> vdd vss nand2
    Xi2 wait_cnt<2> conf_waitcycles<2> waithigh<2> vdd vss nand2
    Xi1 wait_cnt<1> conf_waitcycles<1> waithigh<1> vdd vss nand2
    Xi0 wait_cnt<0> conf_waitcycles<0> waithigh<0> vdd vss nand2
    Xi15 net14 net13 wait_rst_rst' vdd vss nand2
    Xi11 net19 net18 wait_rst vdd vss nand2
    Xi5 wait_rst' rst' cnt_rst vdd vss nand2
    Xi22 net025 net030 net029 vdd vss nor2
    Xi12 edge edge' wait_rst' vdd vss nor2
    Xi6 wait_rst rst cnt_rst' vdd vss nor2
    Xi25 enable_e2l net049 net050 rst rst' vdd vss dff_st_ar_dh
    Xi24 ready wait_ready net034 rst rst' vdd vss dff_st_ar_dh
    Xi8 int edge net18 wait_rst_rst wait_rst_rst' vdd vss dff_st_ar_dh
    Xi7 net15 edge' net19 wait_rst_rst wait_rst_rst' vdd vss dff_st_ar_dh
    Xi23 net029 ready vdd vss inv
    Xi16 wait_rst_rst' wait_rst_rst vdd vss inv
    Xi9 int net15 vdd vss inv
    Xi14 wait_cnt<4> wait_cnt<5> wait_cnt<6> wait_cnt<7> net13 vdd vss nor4
    Xi13 wait_cnt<0> wait_cnt<1> wait_cnt<2> wait_cnt<3> net14 vdd vss nor4
    Xi21 waithigh<0> waithigh<1> waithigh<2> waithigh<3> net025 vdd vss nand4
    Xi20 waithigh<4> waithigh<5> waithigh<6> waithigh<7> net030 vdd vss nand4
    Xi27 net052 clk_int vdd vss buffer
.ENDS

.SUBCKT ff_ready_2 ff0<0> ff0<1> ff1<0> ff1<1> ff_ready rst rst' vdd vss
    Xi2 ff_nor0 ff_nor1 ff_nand vdd vss nand2
    Xi3 ff_nand ff_ready net18 rst rst' vdd vss dff_st_ar_dh
    Xi0 ff0<0> ff0<1> ff_nor0 vdd vss nor2
    Xi1 ff1<0> ff1<1> ff_nor1 vdd vss nor2
.ENDS

.SUBCKT tdc_ready_2 alarm<0> alarm<1> clk conf_maxcycles<0> conf_maxcycles<1> conf_maxcycles<2>
                    + conf_maxcycles<3> conf_maxcycles<4> conf_maxcycles<5> conf_maxcycles<6>
                    + conf_maxcycles<7> conf_waitcycles<0> conf_waitcycles<1> conf_waitcycles<2>
                    + conf_waitcycles<3> conf_waitcycles<4> conf_waitcycles<5> conf_waitcycles<6>
                    + conf_waitcycles<7> enable_e2l ff0<0> ff0<1> ff1<0> ff1<1> int ready rst rst'
                    + vdd vss
    Xi20 conf_maxcycles<0> conf_maxcycles<1> conf_maxcycles<2> conf_maxcycles<3> conf_maxcycles<4>
         + conf_maxcycles<5> conf_maxcycles<6> conf_maxcycles<7> int net017 rst rst' vdd vss
         + max_ready
    Xi32 alarm<0> net19 net027 ready_i vdd vss nand3
    Xi19 clk conf_waitcycles<0> conf_waitcycles<1> conf_waitcycles<2> conf_waitcycles<3>
         + conf_waitcycles<4> conf_waitcycles<5> conf_waitcycles<6> conf_waitcycles<7> enable_e2l
         + int rst rst' vdd vss wait_ready wait_ready
    Xi28 wait_ready net19 vdd vss inv
    Xi27 ff_ready alarm<0> vdd vss inv
    Xi30 ready_i ready ready' rst rst' vdd vss dff_st_ar_dh
    Xi33 net017 ready' alarm<1> net027 rst rst' vdd vss dff_st_ar
    Xi18 ff0<0> ff0<1> ff1<0> ff1<1> ff_ready rst rst' vdd vss ff_ready_2
.ENDS

.SUBCKT tdc_1b_diff_branch alarm<0> alarm<1> buf1_p<0> clk conf0_n<0> conf0_n<1> conf0_n<2>
                           + conf0_n<3> conf0_n<4> conf0_n<5> conf0_n<6> conf0_n<7> conf0_p<0>
                           + conf0_p<1> conf0_p<2> conf0_p<3> conf0_p<4> conf0_p<5> conf0_p<6>
                           + conf0_p<7> conf1_n<0> conf1_n<1> conf1_n<2> conf1_n<3> conf1_n<4>
                           + conf1_n<5> conf1_n<6> conf1_n<7> conf1_p<0> conf1_p<1> conf1_p<2>
                           + conf1_p<3> conf1_p<4> conf1_p<5> conf1_p<6> conf1_p<7> conf_dec<0>
                           + conf_dec<1> conf_dec<2> conf_dec<3> conf_maxcycles<0> conf_maxcycles<1>
                           + conf_maxcycles<2> conf_maxcycles<3> conf_maxcycles<4> conf_maxcycles<5>
                           + conf_maxcycles<6> conf_maxcycles<7> conf_waitcycles<0>
                           + conf_waitcycles<1> conf_waitcycles<2> conf_waitcycles<3>
                           + conf_waitcycles<4> conf_waitcycles<5> conf_waitcycles<6>
                           + conf_waitcycles<7> edge0_n edge0_p edge1_n edge1_p enable_e2l ff<0>
                           + ff<1> ff<2> ff<3> rand_out ready rst rst' vdd vss
    Xi1 net31<0> net31<1> buf0_p<0> buf0_p<1> net30<0> net30<1> buf1_p<0> buf1_p<1> conf0_n<0>
        + conf0_n<1> conf0_n<2> conf0_n<3> conf0_n<4> conf0_n<5> conf0_n<6> conf0_n<7> conf0_p<0>
        + conf0_p<1> conf0_p<2> conf0_p<3> conf0_p<4> conf0_p<5> conf0_p<6> conf0_p<7> conf1_n<0>
        + conf1_n<1> conf1_n<2> conf1_n<3> conf1_n<4> conf1_n<5> conf1_n<6> conf1_n<7> conf1_p<0>
        + conf1_p<1> conf1_p<2> conf1_p<3> conf1_p<4> conf1_p<5> conf1_p<6> conf1_p<7> edge0_n
        + edge0_p edge1_n edge1_p ff<0> ff<1> ff<2> ff<3> rst rst' vdd vss
        + tdc_2e_1b_diff_np_4lin_buf
    Xi7 conf_dec<0> conf_dec<1> conf_dec<2> conf_dec<3> ff<0> ff<1> ff<2> ff<3> rand_out vdd vss
        + dec_4_conf_0
    Xi2 alarm<0> alarm<1> clk conf_maxcycles<0> conf_maxcycles<1> conf_maxcycles<2>
        + conf_maxcycles<3> conf_maxcycles<4> conf_maxcycles<5> conf_maxcycles<6> conf_maxcycles<7>
        + conf_waitcycles<0> conf_waitcycles<1> conf_waitcycles<2> conf_waitcycles<3>
        + conf_waitcycles<4> conf_waitcycles<5> conf_waitcycles<6> conf_waitcycles<7> enable_e2l
        + ff<0> ff<1> ff<2> ff<3> buf0_p<0> ready rst rst' vdd vss tdc_ready_2
.ENDS
