* Top cell name: dc_collection

.SUBCKT buffer in out vdd vss
    Mm1 out int vss vss n_mos l=60n w=480.0n m=4
    Mm0 int in vss vss n_mos l=60n w=480.0n m=1
    Mm3 out int vdd vdd p_mos l=60n w=480.0n m=4
    Mm2 int in vdd vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm5 net17 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm4 net18 in1 net17 vss n_mos l=60n w=360.0n m=1
    Mm3 out in0 net18 vss n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=60n w=360.0n m=1
    Mm2 net5 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm1 net16 in1 net5 vss n_mos l=60n w=360.0n m=1
    Mm0 out in0 net16 vss n_mos l=60n w=360.0n m=1
    Mm7 net32 rst vdd vdd p_mos l=60n w=480.0n m=1
    Mm6 out in2 net32 vdd p_mos l=60n w=480.0n m=1
    Mm5 out in1 net32 vdd p_mos l=60n w=480.0n m=1
    Mm4 out in0 net32 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=120.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT dff_st_ar_buf clk d q q' rst rst' vdd vss
    Xi0 clk d net17 net18 rst rst' vdd vss dff_st_ar
    Xi2 net17 q' vdd vss inv
    Xi1 net18 q vdd vss inv
.ENDS

.SUBCKT edge_to_level_3e edge enable out0 out1 out2 rst rst' vdd vss
    Xi5 edge out1 out2 net17 rst rst' vdd vss dff_st_ar_buf
    Xi4 edge out0 out1 net18 rst rst' vdd vss dff_st_ar_buf
    Xi3 edge enable out0 net19 rst rst' vdd vss dff_st_ar_buf
.ENDS

.SUBCKT mero_nand2 in0 in1 out vdd vss
    Mm1 out in1 vdd vdd p_mos l=60n w=120.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=120.0n m=1
    Mm3 net7 in1 vss vss n_mos l=60n w=120.0n m=1
    Mm2 out in0 net7 vss n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT mero_buf in out vdd vss
    Mm1 out net1 vss vss n_mos l=60n w=120.0n m=1
    Mm0 net1 in vss vss n_mos l=60n w=120.0n m=1
    Mm3 out net1 vdd vdd p_mos l=60n w=120.0n m=1
    Mm2 net1 in vdd vdd p_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT mero_3e_1b enable out0 out1 out2 vdd vss
    Xi2 out1 enable net5 vdd vss mero_nand2
    Xi1 out0 enable net6 vdd vss mero_nand2
    Xi0 out2 enable net7 vdd vss mero_nand2
    Xi5 net5 out2 vdd vss mero_buf
    Xi4 net6 out1 vdd vss mero_buf
    Xi3 net7 out0 vdd vss mero_buf
.ENDS

.SUBCKT nor2 in0 in1 out vdd vss
    Mm1 out in1 vss vss n_mos l=60n w=120.0n m=1
    Mm0 out in0 vss vss n_mos l=60n w=120.0n m=1
    Mm3 net7 in1 vdd vdd p_mos l=60n w=480.0n m=1
    Mm2 out in0 net7 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dc_3e_1b_no_config enable_e2l enable_mero int0 int1 int2 out0 out1 out2 rst rst' vdd vss
    Xi11 mero_out2 int2 vdd vss buffer
    Xi9 mero_out0 int0 vdd vss buffer
    Xi10 mero_out1 int1 vdd vss buffer
    Xi1 int1 enable_e2l out0 out1 out2 rst rst' vdd vss edge_to_level_3e
    Xi5 enable_int mero_out0 mero_out1 mero_out2 vdd vss mero_3e_1b
    Xi12 out2 net10 enable_int vdd vss nor2
    Xi13 enable_mero net10 vdd vss inv
.ENDS

.SUBCKT mero_3e_4b enable out0 out1 out2 vdd vss
    Xi2 out1 enable int2<0> vdd vss mero_nand2
    Xi1 out0 enable int1<0> vdd vss mero_nand2
    Xi0 out2 enable int0<0> vdd vss mero_nand2
    Xi14 int2<3> out2 vdd vss mero_buf
    Xi13 int1<3> out1 vdd vss mero_buf
    Xi12 int0<3> out0 vdd vss mero_buf
    Xi11 int2<2> int2<3> vdd vss mero_buf
    Xi10 int1<2> int1<3> vdd vss mero_buf
    Xi9 int0<2> int0<3> vdd vss mero_buf
    Xi8 int2<1> int2<2> vdd vss mero_buf
    Xi7 int2<0> int2<1> vdd vss mero_buf
    Xi6 int1<1> int1<2> vdd vss mero_buf
    Xi5 int1<0> int1<1> vdd vss mero_buf
    Xi4 int0<1> int0<2> vdd vss mero_buf
    Xi3 int0<0> int0<1> vdd vss mero_buf
.ENDS

.SUBCKT dc_3e_4b_no_config enable_e2l enable_mero int0 int1 int2 out0 out1 out2 rst rst' vdd vss
    Xi11 mero_out2 int2 vdd vss buffer
    Xi9 mero_out0 int0 vdd vss buffer
    Xi10 mero_out1 int1 vdd vss buffer
    Xi1 int1 enable_e2l out0 out1 out2 rst rst' vdd vss edge_to_level_3e
    Xi5 enable_int mero_out0 mero_out1 mero_out2 vdd vss mero_3e_4b
    Xi12 out2 net013 enable_int vdd vss nor2
    Xi13 enable_mero net013 vdd vss inv
.ENDS

.SUBCKT mero_3e_3b enable out0 out1 out2 vdd vss
    Xi2 out1 enable int2<0> vdd vss mero_nand2
    Xi1 out0 enable int1<0> vdd vss mero_nand2
    Xi0 out2 enable int0<0> vdd vss mero_nand2
    Xi14 int2<2> out2 vdd vss mero_buf
    Xi13 int1<2> out1 vdd vss mero_buf
    Xi12 int0<2> out0 vdd vss mero_buf
    Xi8 int2<1> int2<2> vdd vss mero_buf
    Xi7 int2<0> int2<1> vdd vss mero_buf
    Xi6 int1<1> int1<2> vdd vss mero_buf
    Xi5 int1<0> int1<1> vdd vss mero_buf
    Xi4 int0<1> int0<2> vdd vss mero_buf
    Xi3 int0<0> int0<1> vdd vss mero_buf
.ENDS

.SUBCKT dc_3e_3b_no_config enable_e2l enable_mero int0 int1 int2 out0 out1 out2 rst rst' vdd vss
    Xi11 mero_out2 int2 vdd vss buffer
    Xi9 mero_out0 int0 vdd vss buffer
    Xi10 mero_out1 int1 vdd vss buffer
    Xi1 int1 enable_e2l out0 out1 out2 rst rst' vdd vss edge_to_level_3e
    Xi12 out2 net014 enable_int vdd vss nor2
    Xi5 enable_int mero_out0 mero_out1 mero_out2 vdd vss mero_3e_3b
    Xi13 enable_mero net014 vdd vss inv
.ENDS

.SUBCKT single_ended_to_diff in out_n out_p vdd vss
    Mm2 out_n in vdd vdd p_mos l=60n w=480.0n m=4
    Mm3 out_p out_n vdd vdd p_mos l=60n w=480.0n m=4
    Mm1 out_p out_n vss vss n_mos l=60n w=480.0n m=4
    Mm0 out_n in vss vss n_mos l=60n w=480.0n m=4
.ENDS

.SUBCKT mux2 in0 in1 out sel vdd vss
    Xi2 net16 net15 out vdd vss nand2
    Xi1 sel in1 net15 vdd vss nand2
    Xi0 in0 net14 net16 vdd vss nand2
    Mm0 net14 sel vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 net14 sel vss vss n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux4 in<0> in<1> in<2> in<3> out sel<0> sel<1> vdd vss
    Xi2 net8 net7 out sel<1> vdd vss mux2
    Xi1 in<2> in<3> net7 sel<0> vdd vss mux2
    Xi0 in<0> in<1> net8 sel<0> vdd vss mux2
.ENDS

.SUBCKT dec4_inverted out<0> out<1> out<2> out<3> sel<0> sel<1> vdd vss
    Xi1 sel<1> sel'<1> vdd vss inv
    Xi0 sel<0> sel'<0> vdd vss inv
    Xi6 sel<0> sel<1> out<3> vdd vss nand2
    Xi5 sel'<0> sel<1> out<2> vdd vss nand2
    Xi4 sel<0> sel'<1> out<1> vdd vss nand2
    Xi3 sel'<0> sel'<1> out<0> vdd vss nand2
.ENDS

.SUBCKT mero_3e_2b enable out0 out1 out2 vdd vss
    Xi2 out1 enable int2<0> vdd vss mero_nand2
    Xi1 out0 enable int1<0> vdd vss mero_nand2
    Xi0 out2 enable int0<0> vdd vss mero_nand2
    Xi8 int2<1> out2 vdd vss mero_buf
    Xi7 int2<0> int2<1> vdd vss mero_buf
    Xi6 int1<1> out1 vdd vss mero_buf
    Xi5 int1<0> int1<1> vdd vss mero_buf
    Xi4 int0<1> out0 vdd vss mero_buf
    Xi3 int0<0> int0<1> vdd vss mero_buf
.ENDS

.SUBCKT dc_3e_2b_no_config enable_e2l enable_mero int0 int1 int2 out0 out1 out2 rst rst' vdd vss
    Xi5 enable_int mero_out0 mero_out1 mero_out2 vdd vss mero_3e_2b
    Xi1 int1 enable_e2l out0 out1 out2 rst rst' vdd vss edge_to_level_3e
    Xi12 out2 net014 enable_int vdd vss nor2
    Xi9 mero_out0 int0 vdd vss buffer
    Xi11 mero_out2 int2 vdd vss buffer
    Xi10 mero_out1 int1 vdd vss buffer
    Xi13 enable_mero net014 vdd vss inv
.ENDS

.SUBCKT xor2 in0 in1 out vdd vss
    Mm3 out in0' net20 vdd p_mos l=60n w=240.0n m=1
    Mm2 net20 in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in0 net21 vdd p_mos l=60n w=240.0n m=1
    Mm0 net21 in1' vdd vdd p_mos l=60n w=240.0n m=1
    Mm7 net19 in1 vss vss n_mos l=60n w=120.0n m=1
    Mm6 net18 in1' vss vss n_mos l=60n w=120.0n m=1
    Mm5 out in0' net18 vss n_mos l=60n w=120.0n m=1
    Mm4 out in0 net19 vss n_mos l=60n w=120.0n m=1
    Xi1 in1 in1' vdd vss inv
    Xi0 in0 in0' vdd vss inv
.ENDS

.SUBCKT nor3 in0 in1 in2 out vdd vss
    Mm2 out in0 net6 vdd p_mos l=60n w=480.0n m=1
    Mm1 net6 in1 net7 vdd p_mos l=60n w=480.0n m=1
    Mm0 net7 in2 vdd vdd p_mos l=60n w=480.0n m=1
    Mm5 out in2 vss vss n_mos l=60n w=120.0n m=1
    Mm4 out in0 vss vss n_mos l=60n w=120.0n m=1
    Mm3 out in1 vss vss n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT mero_collapse_3e alarm enable_e2l int0 int1 int2 rst rst' vdd vss
    Xi2 int2 int1 xor2 vdd vss xor2
    Xi1 int0 int2 xor1 vdd vss xor2
    Xi0 int1 int0 xor0 vdd vss xor2
    Xi7 nor or vdd vss inv
    Xi4 xor0 xor1 xor2 nor vdd vss nor3
    Xi6 enable_e2l or alarm net016 rst rst' vdd vss dff_st_ar
.ENDS

.SUBCKT vdd_gate_1ma enable' vdd_in vdd_out vss
    Mm0 vdd_out enable' vdd_in vdd_in p_mos_lvt l=60n w=4u m=40
    Mm1 vdd_out enable' vss vss n_mos_lvt l=60n w=4u m=40
.ENDS

.SUBCKT dc_collection alarm_dc conf_seldc<0> conf_seldc<1> dcedge0<1> dcedge0<2> dcedge0<3>
                      + dcedge1<1> dcedge1<2> dcedge1<3> dcedge2<1> dcedge2<2> dcedge2<3> edge0_n
                      + edge0_p edge1_n edge1_p edge2_n edge2_p enable_e2l enable_mero mero_int<0>
                      + mero_int<1> mero_int<2> rst rst' sel_dcedge<0> sel_dcedge<1> vdd_core vdd_dc
                      + vss
    Xi29 enable_e2l enable_mero mero_int0<0> mero_int1<0> mero_int2<0> mero_edge0<0> mero_edge1<0>
         + mero_edge2<0> rst rst' vdd_dc_int<0> vss dc_3e_1b_no_config
    Xi27 enable_e2l enable_mero mero_int0<3> mero_int1<3> mero_int2<3> mero_edge0<3> mero_edge1<3>
         + mero_edge2<3> rst rst' vdd_dc_int<3> vss dc_3e_4b_no_config
    Xi0 enable_e2l enable_mero mero_int0<2> mero_int1<2> mero_int2<2> mero_edge0<2> mero_edge1<2>
        + mero_edge2<2> rst rst' vdd_dc_int<2> vss dc_3e_3b_no_config
    Xi9 sedge0 edge0_n edge0_p vdd_dc vss single_ended_to_diff
    Xi11 sedge1 edge1_n edge1_p vdd_dc vss single_ended_to_diff
    Xi10 sedge2 edge2_n edge2_p vdd_dc vss single_ended_to_diff
    Xi21 mero_edge0<0> mero_edge0<1> mero_edge0<2> mero_edge0<3> dcedge0<0> conf_seldc<0>
         + conf_seldc<1> vdd_core vss mux4
    Xi19 mero_int0<0> mero_int0<1> mero_int0<2> mero_int0<3> mero_int<0> conf_seldc<0> conf_seldc<1>
         + vdd_core vss mux4
    Xi14 dcedge0<0> dcedge0<1> dcedge0<2> dcedge0<3> sedge0 sel_dcedge<0> sel_dcedge<1> vdd_core vss
         + mux4
    Xi22 mero_edge1<0> mero_edge1<1> mero_edge1<2> mero_edge1<3> dcedge1<0> conf_seldc<0>
         + conf_seldc<1> vdd_core vss mux4
    Xi18 mero_int1<0> mero_int1<1> mero_int1<2> mero_int1<3> mero_int<1> conf_seldc<0> conf_seldc<1>
         + vdd_core vss mux4
    Xi15 dcedge1<0> dcedge1<1> dcedge1<2> dcedge1<3> sedge1 sel_dcedge<0> sel_dcedge<1> vdd_core vss
         + mux4
    Xi20 mero_edge2<0> mero_edge2<1> mero_edge2<2> mero_edge2<3> dcedge2<0> conf_seldc<0>
         + conf_seldc<1> vdd_core vss mux4
    Xi17 mero_int2<0> mero_int2<1> mero_int2<2> mero_int2<3> mero_int<2> conf_seldc<0> conf_seldc<1>
         + vdd_core vss mux4
    Xi16 dcedge2<0> dcedge2<1> dcedge2<2> dcedge2<3> sedge2 sel_dcedge<0> sel_dcedge<1> vdd_core vss
         + mux4
    Xi30 seldc_dec<0> seldc_dec<1> seldc_dec<2> seldc_dec<3> conf_seldc<0> conf_seldc<1> vdd_core
         + vss dec4_inverted
    Xi24 enable_e2l enable_mero mero_int0<1> mero_int1<1> mero_int2<1> mero_edge0<1> mero_edge1<1>
         + mero_edge2<1> rst rst' vdd_dc_int<1> vss dc_3e_2b_no_config
    Xi3 alarm_dc enable_e2l mero_int<0> mero_int<1> mero_int<2> rst rst' vdd_dc vss mero_collapse_3e
    Xi28 seldc_dec<0> vdd_dc vdd_dc_int<0> vss vdd_gate_1ma
    Xi26 seldc_dec<3> vdd_dc vdd_dc_int<3> vss vdd_gate_1ma
    Xi25 seldc_dec<1> vdd_dc vdd_dc_int<1> vss vdd_gate_1ma
    Xi23 seldc_dec<2> vdd_dc vdd_dc_int<2> vss vdd_gate_1ma
.ENDS
