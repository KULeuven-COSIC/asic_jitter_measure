* Top cell name: conf_4

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm5 net17 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm4 net18 in1 net17 vss n_mos l=60n w=360.0n m=1
    Mm3 out in0 net18 vss n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=60n w=360.0n m=1
    Mm2 net5 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm1 net16 in1 net5 vss n_mos l=60n w=360.0n m=1
    Mm0 out in0 net16 vss n_mos l=60n w=360.0n m=1
    Mm7 net32 rst vdd vdd p_mos l=60n w=480.0n m=1
    Mm6 out in2 net32 vdd p_mos l=60n w=480.0n m=1
    Mm5 out in1 net32 vdd p_mos l=60n w=480.0n m=1
    Mm4 out in0 net32 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=120.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT dff_st_ar_buf clk d q q' rst rst' vdd vss
    Xi0 clk d net17 net18 rst rst' vdd vss dff_st_ar
    Xi2 net17 q' vdd vss inv
    Xi1 net18 q vdd vss inv
.ENDS

.SUBCKT conf_2 clk in out<0> out<1> rst rst' vdd vss
    Xi1 clk out<0> out<1> net14 rst rst' vdd vss dff_st_ar_buf
    Xi0 clk in out<0> net13 rst rst' vdd vss dff_st_ar_buf
.ENDS

.SUBCKT conf_4 clk in out<0> out<1> out<2> out<3> rst rst' vdd vss
    Xi1 clk out<1> out<2> out<3> rst rst' vdd vss conf_2
    Xi0 clk in out<0> out<1> rst rst' vdd vss conf_2
.ENDS
