* Top cell name: dc_scan_jit_128

.SUBCKT nand2 IN0 IN1 OUT VDD VSS
    Mm1 net13 IN1 VSS VSS n_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 net13 VSS n_mos l=60n w=240.0n m=1
    Mm3 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm2 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 IN0 IN1 IN2 OUT VDD VSS
    Mm2 OUT IN2 VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
    Mm5 net17 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm4 net18 IN1 net17 VSS n_mos l=60n w=360.0n m=1
    Mm3 OUT IN0 net18 VSS n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r IN0 IN1 IN2 OUT RST VDD VSS
    Mm3 OUT RST VSS VSS n_mos l=60n w=360.0n m=1
    Mm2 net5 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm1 net16 IN1 net5 VSS n_mos l=60n w=360.0n m=1
    Mm0 OUT IN0 net16 VSS n_mos l=60n w=360.0n m=1
    Mm7 net32 RST VDD VDD p_mos l=60n w=480.0n m=1
    Mm6 OUT IN2 net32 VDD p_mos l=60n w=480.0n m=1
    Mm5 OUT IN1 net32 VDD p_mos l=60n w=480.0n m=1
    Mm4 OUT IN0 net32 VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar CLK D Q Q' RST RST' VDD VSS
    Xi5 Q N1 Q' VDD VSS nand2
    Xi4 N0 Q' Q VDD VSS nand2
    Xi3 N1 D N3 VDD VSS nand2
    Xi0 N3 N0 N2 VDD VSS nand2
    Xi1 CLK N2 RST' N0 VDD VSS nand3
    Xi2 CLK N0 N3 N1 RST VDD VSS nand3_r
.ENDS

.SUBCKT inv_jit IN OUT VDD VSS
    Mm0 OUT IN VDD VDD p_mos l=60n w=480.0n m=1
    Mm1 OUT IN VSS VSS n_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dc_jit_2 CLK IN LAST OUT<0> OUT<1> RST RST' VDD VSS
    Xi3 CLK LAST OUT<1> net24 RST RST' VDD VSS dff_st_ar
    Xi2 CLK INT net25 OUT<0> RST RST' VDD VSS dff_st_ar
    Xi1 INT LAST VDD VSS inv_jit
    Xi0 IN INT VDD VSS inv_jit
.ENDS

.SUBCKT dc_jit_4 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<2> OUT<3> RST RST' VDD VSS dc_jit_2
    Xi0 CLK IN INT OUT<0> OUT<1> RST RST' VDD VSS dc_jit_2
.ENDS

.SUBCKT dc_jit_8 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD
                 + VSS
    Xi1 CLK INT LAST OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS dc_jit_4
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS dc_jit_4
.ENDS

.SUBCKT dc_jit_16 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS
        + dc_jit_8
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> RST RST' VDD VSS dc_jit_8
.ENDS

.SUBCKT dc_jit_32 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                  + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                  + OUT<30> OUT<31> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25>
        + OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST' VDD VSS dc_jit_16
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> RST RST' VDD VSS dc_jit_16
.ENDS

.SUBCKT dc_jit_64 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                  + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                  + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                  + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                  + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                  + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                  + OUT<60> OUT<61> OUT<62> OUT<63> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41>
        + OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52>
        + OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63>
        + RST RST' VDD VSS dc_jit_32
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21>
        + OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> RST RST'
        + VDD VSS dc_jit_32
.ENDS

.SUBCKT dc_jit_128 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9>
                   + OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19>
                   + OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29>
                   + OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39>
                   + OUT<40> OUT<41> OUT<42> OUT<43> OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49>
                   + OUT<50> OUT<51> OUT<52> OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59>
                   + OUT<60> OUT<61> OUT<62> OUT<63> OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69>
                   + OUT<70> OUT<71> OUT<72> OUT<73> OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79>
                   + OUT<80> OUT<81> OUT<82> OUT<83> OUT<84> OUT<85> OUT<86> OUT<87> OUT<88> OUT<89>
                   + OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95> OUT<96> OUT<97> OUT<98> OUT<99>
                   + OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105> OUT<106> OUT<107>
                   + OUT<108> OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115>
                   + OUT<116> OUT<117> OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123>
                   + OUT<124> OUT<125> OUT<126> OUT<127> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<64> OUT<65> OUT<66> OUT<67> OUT<68> OUT<69> OUT<70> OUT<71> OUT<72> OUT<73>
        + OUT<74> OUT<75> OUT<76> OUT<77> OUT<78> OUT<79> OUT<80> OUT<81> OUT<82> OUT<83> OUT<84>
        + OUT<85> OUT<86> OUT<87> OUT<88> OUT<89> OUT<90> OUT<91> OUT<92> OUT<93> OUT<94> OUT<95>
        + OUT<96> OUT<97> OUT<98> OUT<99> OUT<100> OUT<101> OUT<102> OUT<103> OUT<104> OUT<105>
        + OUT<106> OUT<107> OUT<108> OUT<109> OUT<110> OUT<111> OUT<112> OUT<113> OUT<114> OUT<115>
        + OUT<116> OUT<117> OUT<118> OUT<119> OUT<120> OUT<121> OUT<122> OUT<123> OUT<124> OUT<125>
        + OUT<126> OUT<127> RST RST' VDD VSS dc_jit_64
    Xi0 CLK IN INT OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> OUT<7> OUT<8> OUT<9> OUT<10>
        + OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> OUT<17> OUT<18> OUT<19> OUT<20> OUT<21>
        + OUT<22> OUT<23> OUT<24> OUT<25> OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32>
        + OUT<33> OUT<34> OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43>
        + OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> OUT<53> OUT<54>
        + OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> OUT<62> OUT<63> RST RST' VDD VSS
        + dc_jit_64
.ENDS

.SUBCKT mux2 IN0 IN1 OUT SEL VDD VSS
    Xi2 net16 net15 OUT VDD VSS nand2
    Xi1 SEL IN1 net15 VDD VSS nand2
    Xi0 IN0 net14 net16 VDD VSS nand2
    Mm0 net14 SEL VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 net14 SEL VSS VSS n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT scan_jit_2 CLK IN_PAR<0> IN_PAR<1> IN_SER OUT RST RST' SER VDD VSS
    Xi1 CLK net12 OUT net14 RST RST' VDD VSS dff_st_ar
    Xi0 CLK net07 net11 net15 RST RST' VDD VSS dff_st_ar
    Xi4 IN_PAR<0> IN_SER net07 SER VDD VSS mux2
    Xi2 IN_PAR<1> net11 net12 SER VDD VSS mux2
.ENDS

.SUBCKT scan_jit_4 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_SER net8 RST RST' SER VDD VSS scan_jit_2
    Xi6 CLK IN_PAR<2> IN_PAR<3> net8 OUT RST RST' SER VDD VSS scan_jit_2
.ENDS

.SUBCKT scan_jit_8 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                   + IN_PAR<7> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_SER net8 RST RST' SER VDD VSS scan_jit_4
    Xi6 CLK IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> net8 OUT RST RST' SER VDD VSS scan_jit_4
.ENDS

.SUBCKT scan_jit_16 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7> IN_SER
        + net8 RST RST' SER VDD VSS scan_jit_8
    Xi6 CLK IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + net8 OUT RST RST' SER VDD VSS scan_jit_8
.ENDS

.SUBCKT scan_jit_32 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                    + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                    + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_16
    Xi6 CLK IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + net8 OUT RST RST' SER VDD VSS scan_jit_16
.ENDS

.SUBCKT scan_jit_64 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                    + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                    + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                    + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                    + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_PAR<32> IN_PAR<33> IN_PAR<34>
                    + IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39> IN_PAR<40> IN_PAR<41>
                    + IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47> IN_PAR<48>
                    + IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
                    + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62>
                    + IN_PAR<63> IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_32
    Xi6 CLK IN_PAR<32> IN_PAR<33> IN_PAR<34> IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39>
        + IN_PAR<40> IN_PAR<41> IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47>
        + IN_PAR<48> IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
        + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62> IN_PAR<63>
        + net8 OUT RST RST' SER VDD VSS scan_jit_32
.ENDS

.SUBCKT scan_jit_128 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6>
                     + IN_PAR<7> IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13>
                     + IN_PAR<14> IN_PAR<15> IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20>
                     + IN_PAR<21> IN_PAR<22> IN_PAR<23> IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27>
                     + IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31> IN_PAR<32> IN_PAR<33> IN_PAR<34>
                     + IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39> IN_PAR<40> IN_PAR<41>
                     + IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47> IN_PAR<48>
                     + IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
                     + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62>
                     + IN_PAR<63> IN_PAR<64> IN_PAR<65> IN_PAR<66> IN_PAR<67> IN_PAR<68> IN_PAR<69>
                     + IN_PAR<70> IN_PAR<71> IN_PAR<72> IN_PAR<73> IN_PAR<74> IN_PAR<75> IN_PAR<76>
                     + IN_PAR<77> IN_PAR<78> IN_PAR<79> IN_PAR<80> IN_PAR<81> IN_PAR<82> IN_PAR<83>
                     + IN_PAR<84> IN_PAR<85> IN_PAR<86> IN_PAR<87> IN_PAR<88> IN_PAR<89> IN_PAR<90>
                     + IN_PAR<91> IN_PAR<92> IN_PAR<93> IN_PAR<94> IN_PAR<95> IN_PAR<96> IN_PAR<97>
                     + IN_PAR<98> IN_PAR<99> IN_PAR<100> IN_PAR<101> IN_PAR<102> IN_PAR<103>
                     + IN_PAR<104> IN_PAR<105> IN_PAR<106> IN_PAR<107> IN_PAR<108> IN_PAR<109>
                     + IN_PAR<110> IN_PAR<111> IN_PAR<112> IN_PAR<113> IN_PAR<114> IN_PAR<115>
                     + IN_PAR<116> IN_PAR<117> IN_PAR<118> IN_PAR<119> IN_PAR<120> IN_PAR<121>
                     + IN_PAR<122> IN_PAR<123> IN_PAR<124> IN_PAR<125> IN_PAR<126> IN_PAR<127>
                     + IN_SER OUT RST RST' SER VDD VSS
    Xi5 CLK IN_PAR<0> IN_PAR<1> IN_PAR<2> IN_PAR<3> IN_PAR<4> IN_PAR<5> IN_PAR<6> IN_PAR<7>
        + IN_PAR<8> IN_PAR<9> IN_PAR<10> IN_PAR<11> IN_PAR<12> IN_PAR<13> IN_PAR<14> IN_PAR<15>
        + IN_PAR<16> IN_PAR<17> IN_PAR<18> IN_PAR<19> IN_PAR<20> IN_PAR<21> IN_PAR<22> IN_PAR<23>
        + IN_PAR<24> IN_PAR<25> IN_PAR<26> IN_PAR<27> IN_PAR<28> IN_PAR<29> IN_PAR<30> IN_PAR<31>
        + IN_PAR<32> IN_PAR<33> IN_PAR<34> IN_PAR<35> IN_PAR<36> IN_PAR<37> IN_PAR<38> IN_PAR<39>
        + IN_PAR<40> IN_PAR<41> IN_PAR<42> IN_PAR<43> IN_PAR<44> IN_PAR<45> IN_PAR<46> IN_PAR<47>
        + IN_PAR<48> IN_PAR<49> IN_PAR<50> IN_PAR<51> IN_PAR<52> IN_PAR<53> IN_PAR<54> IN_PAR<55>
        + IN_PAR<56> IN_PAR<57> IN_PAR<58> IN_PAR<59> IN_PAR<60> IN_PAR<61> IN_PAR<62> IN_PAR<63>
        + IN_SER net8 RST RST' SER VDD VSS scan_jit_64
    Xi6 CLK IN_PAR<64> IN_PAR<65> IN_PAR<66> IN_PAR<67> IN_PAR<68> IN_PAR<69> IN_PAR<70> IN_PAR<71>
        + IN_PAR<72> IN_PAR<73> IN_PAR<74> IN_PAR<75> IN_PAR<76> IN_PAR<77> IN_PAR<78> IN_PAR<79>
        + IN_PAR<80> IN_PAR<81> IN_PAR<82> IN_PAR<83> IN_PAR<84> IN_PAR<85> IN_PAR<86> IN_PAR<87>
        + IN_PAR<88> IN_PAR<89> IN_PAR<90> IN_PAR<91> IN_PAR<92> IN_PAR<93> IN_PAR<94> IN_PAR<95>
        + IN_PAR<96> IN_PAR<97> IN_PAR<98> IN_PAR<99> IN_PAR<100> IN_PAR<101> IN_PAR<102>
        + IN_PAR<103> IN_PAR<104> IN_PAR<105> IN_PAR<106> IN_PAR<107> IN_PAR<108> IN_PAR<109>
        + IN_PAR<110> IN_PAR<111> IN_PAR<112> IN_PAR<113> IN_PAR<114> IN_PAR<115> IN_PAR<116>
        + IN_PAR<117> IN_PAR<118> IN_PAR<119> IN_PAR<120> IN_PAR<121> IN_PAR<122> IN_PAR<123>
        + IN_PAR<124> IN_PAR<125> IN_PAR<126> IN_PAR<127> net8 OUT RST RST' SER VDD VSS scan_jit_64
.ENDS

.SUBCKT dc_scan_jit_128 DC_CLK DC_IN DC_LAST DC_RST DC_RST' SCAN_CLK SCAN_IN_SER SCAN_OUT SCAN_RST
                        + SCAN_RST' SCAN_SER VDD VSS
    Xi0 DC_CLK DC_IN DC_LAST DC_OUT<0> DC_OUT<1> DC_OUT<2> DC_OUT<3> DC_OUT<4> DC_OUT<5> DC_OUT<6>
        + DC_OUT<7> DC_OUT<8> DC_OUT<9> DC_OUT<10> DC_OUT<11> DC_OUT<12> DC_OUT<13> DC_OUT<14>
        + DC_OUT<15> DC_OUT<16> DC_OUT<17> DC_OUT<18> DC_OUT<19> DC_OUT<20> DC_OUT<21> DC_OUT<22>
        + DC_OUT<23> DC_OUT<24> DC_OUT<25> DC_OUT<26> DC_OUT<27> DC_OUT<28> DC_OUT<29> DC_OUT<30>
        + DC_OUT<31> DC_OUT<32> DC_OUT<33> DC_OUT<34> DC_OUT<35> DC_OUT<36> DC_OUT<37> DC_OUT<38>
        + DC_OUT<39> DC_OUT<40> DC_OUT<41> DC_OUT<42> DC_OUT<43> DC_OUT<44> DC_OUT<45> DC_OUT<46>
        + DC_OUT<47> DC_OUT<48> DC_OUT<49> DC_OUT<50> DC_OUT<51> DC_OUT<52> DC_OUT<53> DC_OUT<54>
        + DC_OUT<55> DC_OUT<56> DC_OUT<57> DC_OUT<58> DC_OUT<59> DC_OUT<60> DC_OUT<61> DC_OUT<62>
        + DC_OUT<63> DC_OUT<64> DC_OUT<65> DC_OUT<66> DC_OUT<67> DC_OUT<68> DC_OUT<69> DC_OUT<70>
        + DC_OUT<71> DC_OUT<72> DC_OUT<73> DC_OUT<74> DC_OUT<75> DC_OUT<76> DC_OUT<77> DC_OUT<78>
        + DC_OUT<79> DC_OUT<80> DC_OUT<81> DC_OUT<82> DC_OUT<83> DC_OUT<84> DC_OUT<85> DC_OUT<86>
        + DC_OUT<87> DC_OUT<88> DC_OUT<89> DC_OUT<90> DC_OUT<91> DC_OUT<92> DC_OUT<93> DC_OUT<94>
        + DC_OUT<95> DC_OUT<96> DC_OUT<97> DC_OUT<98> DC_OUT<99> DC_OUT<100> DC_OUT<101> DC_OUT<102>
        + DC_OUT<103> DC_OUT<104> DC_OUT<105> DC_OUT<106> DC_OUT<107> DC_OUT<108> DC_OUT<109>
        + DC_OUT<110> DC_OUT<111> DC_OUT<112> DC_OUT<113> DC_OUT<114> DC_OUT<115> DC_OUT<116>
        + DC_OUT<117> DC_OUT<118> DC_OUT<119> DC_OUT<120> DC_OUT<121> DC_OUT<122> DC_OUT<123>
        + DC_OUT<124> DC_OUT<125> DC_OUT<126> DC_OUT<127> DC_RST DC_RST' VDD VSS dc_jit_128
    Xi1 SCAN_CLK DC_OUT<0> DC_OUT<1> DC_OUT<2> DC_OUT<3> DC_OUT<4> DC_OUT<5> DC_OUT<6> DC_OUT<7>
        + DC_OUT<8> DC_OUT<9> DC_OUT<10> DC_OUT<11> DC_OUT<12> DC_OUT<13> DC_OUT<14> DC_OUT<15>
        + DC_OUT<16> DC_OUT<17> DC_OUT<18> DC_OUT<19> DC_OUT<20> DC_OUT<21> DC_OUT<22> DC_OUT<23>
        + DC_OUT<24> DC_OUT<25> DC_OUT<26> DC_OUT<27> DC_OUT<28> DC_OUT<29> DC_OUT<30> DC_OUT<31>
        + DC_OUT<32> DC_OUT<33> DC_OUT<34> DC_OUT<35> DC_OUT<36> DC_OUT<37> DC_OUT<38> DC_OUT<39>
        + DC_OUT<40> DC_OUT<41> DC_OUT<42> DC_OUT<43> DC_OUT<44> DC_OUT<45> DC_OUT<46> DC_OUT<47>
        + DC_OUT<48> DC_OUT<49> DC_OUT<50> DC_OUT<51> DC_OUT<52> DC_OUT<53> DC_OUT<54> DC_OUT<55>
        + DC_OUT<56> DC_OUT<57> DC_OUT<58> DC_OUT<59> DC_OUT<60> DC_OUT<61> DC_OUT<62> DC_OUT<63>
        + DC_OUT<64> DC_OUT<65> DC_OUT<66> DC_OUT<67> DC_OUT<68> DC_OUT<69> DC_OUT<70> DC_OUT<71>
        + DC_OUT<72> DC_OUT<73> DC_OUT<74> DC_OUT<75> DC_OUT<76> DC_OUT<77> DC_OUT<78> DC_OUT<79>
        + DC_OUT<80> DC_OUT<81> DC_OUT<82> DC_OUT<83> DC_OUT<84> DC_OUT<85> DC_OUT<86> DC_OUT<87>
        + DC_OUT<88> DC_OUT<89> DC_OUT<90> DC_OUT<91> DC_OUT<92> DC_OUT<93> DC_OUT<94> DC_OUT<95>
        + DC_OUT<96> DC_OUT<97> DC_OUT<98> DC_OUT<99> DC_OUT<100> DC_OUT<101> DC_OUT<102>
        + DC_OUT<103> DC_OUT<104> DC_OUT<105> DC_OUT<106> DC_OUT<107> DC_OUT<108> DC_OUT<109>
        + DC_OUT<110> DC_OUT<111> DC_OUT<112> DC_OUT<113> DC_OUT<114> DC_OUT<115> DC_OUT<116>
        + DC_OUT<117> DC_OUT<118> DC_OUT<119> DC_OUT<120> DC_OUT<121> DC_OUT<122> DC_OUT<123>
        + DC_OUT<124> DC_OUT<125> DC_OUT<126> DC_OUT<127> SCAN_IN_SER SCAN_OUT SCAN_RST SCAN_RST'
        + SCAN_SER VDD VSS scan_jit_128
.ENDS
