* Top cell name: mux2_10x

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux2 in0 in1 out sel vdd vss
    Xi2 net16 net15 out vdd vss nand2
    Xi1 sel in1 net15 vdd vss nand2
    Xi0 in0 net14 net16 vdd vss nand2
    Mm0 net14 sel vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 net14 sel vss vss n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux2_10x in0<0> in0<1> in0<2> in0<3> in0<4> in0<5> in0<6> in0<7> in0<8> in0<9> in1<0> in1<1>
                 + in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> in1<9> out<0> out<1> out<2>
                 + out<3> out<4> out<5> out<6> out<7> out<8> out<9> sel vdd vss
    Xi0 in0<0> in1<0> out<0> sel vdd vss mux2
    Xi9 in0<9> in1<9> out<9> sel vdd vss mux2
    Xi8 in0<8> in1<8> out<8> sel vdd vss mux2
    Xi7 in0<7> in1<7> out<7> sel vdd vss mux2
    Xi6 in0<6> in1<6> out<6> sel vdd vss mux2
    Xi5 in0<5> in1<5> out<5> sel vdd vss mux2
    Xi4 in0<4> in1<4> out<4> sel vdd vss mux2
    Xi3 in0<3> in1<3> out<3> sel vdd vss mux2
    Xi2 in0<2> in1<2> out<2> sel vdd vss mux2
    Xi1 in0<1> in1<1> out<1> sel vdd vss mux2
.ENDS
