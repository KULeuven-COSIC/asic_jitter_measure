* Top cell name: dc_jit_4

.SUBCKT nand2 IN0 IN1 OUT VDD VSS
    Mm1 net13 IN1 VSS VSS n_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 net13 VSS n_mos l=60n w=240.0n m=1
    Mm3 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm2 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT nand3 IN0 IN1 IN2 OUT VDD VSS
    Mm2 OUT IN2 VDD VDD p_mos l=60n w=240.0n m=1
    Mm1 OUT IN1 VDD VDD p_mos l=60n w=240.0n m=1
    Mm0 OUT IN0 VDD VDD p_mos l=60n w=240.0n m=1
    Mm5 net17 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm4 net18 IN1 net17 VSS n_mos l=60n w=360.0n m=1
    Mm3 OUT IN0 net18 VSS n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r IN0 IN1 IN2 OUT RST VDD VSS
    Mm3 OUT RST VSS VSS n_mos l=60n w=360.0n m=1
    Mm2 net5 IN2 VSS VSS n_mos l=60n w=360.0n m=1
    Mm1 net16 IN1 net5 VSS n_mos l=60n w=360.0n m=1
    Mm0 OUT IN0 net16 VSS n_mos l=60n w=360.0n m=1
    Mm7 net32 RST VDD VDD p_mos l=60n w=480.0n m=1
    Mm6 OUT IN2 net32 VDD p_mos l=60n w=480.0n m=1
    Mm5 OUT IN1 net32 VDD p_mos l=60n w=480.0n m=1
    Mm4 OUT IN0 net32 VDD p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar CLK D Q Q' RST RST' VDD VSS
    Xi5 Q N1 Q' VDD VSS nand2
    Xi4 N0 Q' Q VDD VSS nand2
    Xi3 N1 D N3 VDD VSS nand2
    Xi0 N3 N0 N2 VDD VSS nand2
    Xi1 CLK N2 RST' N0 VDD VSS nand3
    Xi2 CLK N0 N3 N1 RST VDD VSS nand3_r
.ENDS

.SUBCKT inv_jit IN OUT VDD VSS
    Mm0 OUT IN VDD VDD p_mos l=60n w=480.0n m=1
    Mm1 OUT IN VSS VSS n_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dc_jit_2 CLK IN LAST OUT<0> OUT<1> RST RST' VDD VSS
    Xi3 CLK LAST OUT<1> net24 RST RST' VDD VSS dff_st_ar
    Xi2 CLK INT net25 OUT<0> RST RST' VDD VSS dff_st_ar
    Xi1 INT LAST VDD VSS inv_jit
    Xi0 IN INT VDD VSS inv_jit
.ENDS

.SUBCKT dc_jit_4 CLK IN LAST OUT<0> OUT<1> OUT<2> OUT<3> RST RST' VDD VSS
    Xi1 CLK INT LAST OUT<2> OUT<3> RST RST' VDD VSS dc_jit_2
    Xi0 CLK IN INT OUT<0> OUT<1> RST RST' VDD VSS dc_jit_2
.ENDS
