* Top cell name: cal_tdc

.SUBCKT inv_conf conf'<0> conf'<1> conf'<2> conf'<3> conf<0> conf<1> conf<2> conf<3> in out vdd vss
    Mm16 out in vdd vdd p_mos l=60n w=120.0n m=1
    Mm7 out in net16 vdd p_mos l=60n w=120.0n m=1
    Mm6 out in net17 vdd p_mos l=60n w=120.0n m=1
    Mm5 out in net18 vdd p_mos l=60n w=120.0n m=1
    Mm4 out in net19 vdd p_mos l=60n w=120.0n m=1
    Mm3 net16 conf'<3> vdd vdd p_mos l=60n w=120.0n m=1
    Mm2 net17 conf'<2> vdd vdd p_mos l=60n w=120.0n m=1
    Mm1 net18 conf'<1> vdd vdd p_mos l=60n w=120.0n m=1
    Mm0 net19 conf'<0> vdd vdd p_mos l=60n w=120.0n m=1
    Mm17 out in vss vss n_mos l=60n w=120.0n m=1
    Mm15 net20 conf<3> vss vss n_mos l=60n w=120.0n m=1
    Mm14 out in net20 vss n_mos l=60n w=120.0n m=1
    Mm13 net21 conf<2> vss vss n_mos l=60n w=120.0n m=1
    Mm12 out in net21 vss n_mos l=60n w=120.0n m=1
    Mm11 net22 conf<1> vss vss n_mos l=60n w=120.0n m=1
    Mm10 out in net22 vss n_mos l=60n w=120.0n m=1
    Mm9 net23 conf<0> vss vss n_mos l=60n w=120.0n m=1
    Mm8 out in net23 vss n_mos l=60n w=120.0n m=1
.ENDS

.SUBCKT nand2 in0 in1 out vdd vss
    Mm1 net13 in1 vss vss n_mos l=60n w=240.0n m=1
    Mm0 out in0 net13 vss n_mos l=60n w=240.0n m=1
    Mm3 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm2 out in0 vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT ro_2i conf'<0> conf'<1> conf'<2> conf'<3> conf'<4> conf'<5> conf'<6> conf'<7> conf<0>
              + conf<1> conf<2> conf<3> conf<4> conf<5> conf<6> conf<7> enable out vdd vss
    Xi1 conf'<4> conf'<5> conf'<6> conf'<7> conf<4> conf<5> conf<6> conf<7> int out vdd vss inv_conf
    Xi0 conf'<0> conf'<1> conf'<2> conf'<3> conf<0> conf<1> conf<2> conf<3> nand_out int vdd vss
        + inv_conf
    Xi2 out enable nand_out vdd vss nand2
.ENDS

.SUBCKT nand3 in0 in1 in2 out vdd vss
    Mm2 out in2 vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 out in1 vdd vdd p_mos l=60n w=240.0n m=1
    Mm0 out in0 vdd vdd p_mos l=60n w=240.0n m=1
    Mm5 net17 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm4 net18 in1 net17 vss n_mos l=60n w=360.0n m=1
    Mm3 out in0 net18 vss n_mos l=60n w=360.0n m=1
.ENDS

.SUBCKT nand3_r in0 in1 in2 out rst vdd vss
    Mm3 out rst vss vss n_mos l=60n w=360.0n m=1
    Mm2 net5 in2 vss vss n_mos l=60n w=360.0n m=1
    Mm1 net16 in1 net5 vss n_mos l=60n w=360.0n m=1
    Mm0 out in0 net16 vss n_mos l=60n w=360.0n m=1
    Mm7 net32 rst vdd vdd p_mos l=60n w=480.0n m=1
    Mm6 out in2 net32 vdd p_mos l=60n w=480.0n m=1
    Mm5 out in1 net32 vdd p_mos l=60n w=480.0n m=1
    Mm4 out in0 net32 vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT dff_st_ar clk d q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi3 n1 d n3 vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
.ENDS

.SUBCKT tff_st_ar clk q q' rst rst' vdd vss
    Xi0 clk q' q q' rst rst' vdd vss dff_st_ar
.ENDS

.SUBCKT freqscaler3 clk out<0> out<1> out<2> rst rst' vdd vss
    Xi2 int<1> out<2> net16 rst rst' vdd vss tff_st_ar
    Xi1 int<0> out<1> int<1> rst rst' vdd vss tff_st_ar
    Xi0 clk out<0> int<0> rst rst' vdd vss tff_st_ar
.ENDS

.SUBCKT inv_sd in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=480.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT mux2 in0 in1 out sel vdd vss
    Xi2 net16 net15 out vdd vss nand2
    Xi1 sel in1 net15 vdd vss nand2
    Xi0 in0 net14 net16 vdd vss nand2
    Mm0 net14 sel vdd vdd p_mos l=60n w=240.0n m=1
    Mm1 net14 sel vss vss n_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT mux4 in<0> in<1> in<2> in<3> out sel<0> sel<1> vdd vss
    Xi2 net8 net7 out sel<1> vdd vss mux2
    Xi1 in<2> in<3> net7 sel<0> vdd vss mux2
    Xi0 in<0> in<1> net8 sel<0> vdd vss mux2
.ENDS

.SUBCKT inv in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=120.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT inv_bank_8 in<0> in<1> in<2> in<3> in<4> in<5> in<6> in<7> out<0> out<1> out<2> out<3>
                   + out<4> out<5> out<6> out<7> vdd vss
    Xi7 in<7> out<7> vdd vss inv
    Xi6 in<6> out<6> vdd vss inv
    Xi5 in<5> out<5> vdd vss inv
    Xi4 in<4> out<4> vdd vss inv
    Xi3 in<3> out<3> vdd vss inv
    Xi2 in<2> out<2> vdd vss inv
    Xi1 in<1> out<1> vdd vss inv
    Xi0 in<0> out<0> vdd vss inv
.ENDS

.SUBCKT inv_wn in out vdd vss
    Mm0 out in vss vss n_mos l=60n w=240.0n m=1
    Mm1 out in vdd vdd p_mos l=60n w=240.0n m=1
.ENDS

.SUBCKT dff_st_ar_dh clk q q' rst rst' vdd vss
    Xi5 q n1 q' vdd vss nand2
    Xi4 n0 q' q vdd vss nand2
    Xi0 n3 n0 n2 vdd vss nand2
    Xi1 clk n2 rst' n0 vdd vss nand3
    Xi2 clk n0 n3 n1 rst vdd vss nand3_r
    Xi6 n1 n3 vdd vss inv_wn
.ENDS

.SUBCKT dff_st_ar_buf clk d q q' rst rst' vdd vss
    Xi0 clk d net17 net18 rst rst' vdd vss dff_st_ar
    Xi2 net17 q' vdd vss inv
    Xi1 net18 q vdd vss inv
.ENDS

.SUBCKT buffer in out vdd vss
    Mm1 out int vss vss n_mos l=60n w=480.0n m=4
    Mm0 int in vss vss n_mos l=60n w=480.0n m=1
    Mm3 out int vdd vdd p_mos l=60n w=480.0n m=4
    Mm2 int in vdd vdd p_mos l=60n w=480.0n m=1
.ENDS

.SUBCKT cal_tdc cal_enable conf<0> conf<1> conf<2> conf<3> conf<4> conf<5> conf<6> conf<7> out0 out1
                + out2 ro_enable ro_out rst rst' sel<0> sel<1> vdd vss
    Xi0 net6<0> net6<1> net6<2> net6<3> net6<4> net6<5> net6<6> net6<7> conf<0> conf<1> conf<2>
        + conf<3> conf<4> conf<5> conf<6> conf<7> ro_enable ro<0> vdd vss ro_2i
    Xi1 ro<0> ro<1> ro<2> ro<3> rst rst' vdd vss freqscaler3
    Xi8 net023 out0_i vdd vss inv_sd
    Xi4 ro<0> ro<1> ro<2> ro<3> mux_out sel<0> sel<1> vdd vss mux4
    Xi5 conf<0> conf<1> conf<2> conf<3> conf<4> conf<5> conf<6> conf<7> net6<0> net6<1> net6<2>
        + net6<3> net6<4> net6<5> net6<6> net6<7> vdd vss inv_bank_8
    Xi7 cal_enable net027 net023 rst rst' vdd vss dff_st_ar_dh
    Xi3 ro_out out1_i out2_i net11 rst rst' vdd vss dff_st_ar_buf
    Xi2 ro_out cal_enable out1_i net17 rst rst' vdd vss dff_st_ar_buf
    Xi12 out2_i out2 vdd vss buffer
    Xi11 out1_i out1 vdd vss buffer
    Xi10 out0_i out0 vdd vss buffer
    Xi9 mux_out ro_out vdd vss buffer
.ENDS
